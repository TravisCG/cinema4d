MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���om��om��om�}!���om����om��ǔ�om�����om��ol��om��Ɣ�om�����om����om�Rich�om�                        PE  L 1�Q        � !
     �      @-                             0    �  @                   � K   t� (    � �                   � x                                  �� @                                        .text   ��                         `.rdata  ;�     �                @  @.data   �5   �     �             @  �.rsrc   �   �     �             @  @.reloc  N>   �  @   �             @  B                                                                                                                                                                                                                                                                                                                                                U����   SVWQ������9   ������Y�M�j hp�� ����;   �� ���P�o  ���� ����   �   _^[���   ;��<  ��]� ������U����   SVWQ��4����3   ������Y�M���E�P� ��Q�B�Ѓ�;���  ��EPj��MQ�U�R� ��H�Q�҃�;���  �E�_^[���   ;��  ��]� ���������������U����   SVWQ��4����3   ������Y�M���E�P� ��Q�B�Ѓ�;��_  _^[���   ;��O  ��]������������U���0  SVW�������L   ������h�� ���PhD�j�  �������������� t�������  �������
ǅ����    j h����������j h���,�������������Qj h��������l���P�����R������  ���r   Pj ��,���PhJ ��  ��������������  ������������,����������������������_^[��0  ;��#  ��]����������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]��U����   SVWQ��4����3   ������Y�M��M��   �E�� ��E�_^[���   ;��  ��]������U����   SVWQ��4����3   ������Y�M��M��   �E��t�E�P��  ���E�_^[���   ;��>  ��]� ��������U����   SVWQ��4����3   ������Y�M��M��	  �E��  �E�_^[���   ;���  ��]������U����   SVWQ��4����3   ������Y�M��M��   _^[���   ;��  ��]��U����   SVWQ��4����3   ������Y�M��M��	  _^[���   ;��e  ��]��U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�  ���E�_^[���   ;��  ��]� ��������U����   SVW��@����0   ������������u3���   _^[���   ;���  ��]�������������U����   SVW��@����0   ������_^[��]������������U����   SVW��@����0   ������3�_^[��]����������U����   SVWQ��4����3   ������Y�M���E�P� ��Q�B�Ѓ�;��  �E�_^[���   ;���  ��]���������U����   SVW��@����0   ������j0j �)   ��P�EP��  ��_^[���   ;��  ��]������U����   SVW��@����0   ������EE_^[��]������U����   SVW��@����0   ������E� �� �� _^[��]�������������U����   SVW��@����0   ������EP�M���   Q�UR��  ��_^[���   ;���  ��]�����U���  SVWQ��\����i   ������Y�M��X  �M���E��8 u��   �EP��l�����  j h`�������U���P��������  j j���l���Q������R������P�  ��P������Q��
  ��P�����R��
  ��P�E���}  ������؈�c���������	  �������x	  �������m	  �������b	  �������G�����l����L	  ��c�����t�E�P�  ���E�_^[�Ĥ  ;��  ��]� ������������U����   SVWQ��4����3   ������Y�M��E�P�d  ��_^[���   ;��a  ��]��������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��M������E_^[���   ;��  ��]� ������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ��U����   SVWQ��4����3   ������Y�M�3�_^[��]� ��U���  SVW��x����b   ������} u3��   j h�   ��<���P�2������E��\����E��|����E�E��E��<���ǅ@���  �E�  �E�  �E�P �E� �E�p �E�0 �E�@ �E�` h�   ��<���P�MQ�URj�a  ��R��P�� ��  XZ_^[�Ĉ  ;��  ��]Ð   � <����   � np ̋�`����������̋�` ����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`�����������U����   SVW��4����3   ������}s�E   �E��P�i  ���E��}� u3��:�} t�E��Pj �M�Q��  ���E�� �����E����E��$�   �E�_^[���   ;��  ��]������������U����   SVW��4����3   ������} tF�E�E��=$� t�E�x��u�E��P��  �����E�P� ��Q��Ѓ�;��  _^[���   ;��  ��]���U����   SVW��<����1   ������= � tI�}sǅ<���   �	�E��<�����MQ�UR��<���P� ��Q���   �Ѓ�;��  �j�EP�e�����_^[���   ;��r  ��]���������������U����   SVWQ��4����3   ������Y�M��E�� h�E�_^[��]�����������U����   SVWQ��4����3   ������Y�M��M��5   �E��t�E�P�d������E�_^[���   ;���  ��]� ��������U����   SVWQ��4����3   ������Y�M��E�� h_^[��]��������������U����   SVWQ������=   ������Y�M��E��E�}� tM�E쉅 ����� ������������� t%��j��������������;��  ������
ǅ���    �E�    _^[���   ;���
  ��]����������U����   SVW��@����0   �������EP�MQ� ��B�H@�у�;��
  _^[���   ;��
  ��]�������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�.  � ��B���   �у�;��,
  _^[���   ;��
  ��]���������U����   SVWQ��4����3   ������Y�M��M�������E�P� ��Q$�BD�Ѓ�;���	  �E�_^[���   ;��	  ��]�U����   SVWQ��4����3   ������Y�M��M��5�����E�P� ��Q$�BD�Ѓ�;��g	  ��EP�M�Q� ��B$�H�у�;��E	  �E�_^[���   ;��2	  ��]� ������������U����   SVWQ��4����3   ������Y�M��M�������E�P� ��Q$�BD�Ѓ�;���  ��E�P�MQ� ��B$�HL�у�;��  �E�_^[���   ;��  ��]� ������������U����   SVWQ��4����3   ������Y�M���E�P� ��Q$�BH�Ѓ�;��O  �M�����_^[���   ;��7  ��]����U����   SVWQ������<   ������Y�M���E�P�����Q� ��B$�H �у�;���  P�M����������D����E_^[���   ;���  ��]� �����������U����   SVWQ��4����3   ������Y�M���E�P�MQ� ��B$�HL�у�;��k  �E�_^[���   ;��X  ��]� ��U����   SVW������9   ������EP�M�������EP�M�Q� ��B$�H@�у�;��  �E�P�M������M��`����ER��P��" �  XZ_^[���   ;���  ��]�   �" ����   �" fn �U���$  SVW�������I   ������ǅ8���    �= � t!������P� ��=�����8����������������C�����8���������������������������R�M������8�����t��8����������~�����8�����t��8�����������a����E_^[��$  ;���  ��]�����������U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� �����U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�������������U����   SVWQ��4����3   ������Y�M��M��   _^[���   ;���  ��]��U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q� ��B<�H�у�;��  �E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� ����>   ������
ǅ���    �E��@    _^[���   ;��  ��]���������������U����   SVWQ��4����3   ������Y�M��M��E����E��t�E�P�D������E�_^[���   ;��  ��]� ��������U����   SVW��@����0   ������(�����_^[���   ;��h  ��]�����U����   SVW��@����0   ������ ��H����;��-  _^[���   ;��  ��]����������U����   SVW��@����0   �������E�Q� ��B�H�у�;���  �E�     _^[���   ;��  ��]������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P� ��Q�B�Ѓ�;��c  _^[���   ;��S  ��]� �������������U����   SVW��<����1   ������E��<�����<���t��E�(��E�$��   _^[��]� U����   SVW������:   ������E�����������������������q  ������$�|) �   �]  �,����,��=,���   �EP������=�.  }
������&  �} u
������  hp�P���PhD�j�5������� ����� ��� t�� �������������
ǅ���    ������ ��= � t�EP� ��2����   �   �EP�MQ�K�������u����   �   �|�����u�,����,�u\�����������= � t?� ���8�����8�����,�����,��� tj��,����_���������
ǅ���    � �    �   ����_^[���   ;��)   ��]Ð
( �( �(  ( d) �( ������������u�U��� PRSVW�Ej P�w  ��_^[ZX��]�����������̋�U��QSVW3���ى}�9>~H���$    ��F�8�|�����u�T8с<����t�L8�UQR��  ���E�@���E�;|�_^[��]�����������̀=E� uj jj j j �E���  P�{  ����������jjj j j �  ���������������̋�U��Q�M��E�� ��M�Q�  ����]��������������̋�U��Q�M��M������E��t�M�Q�>������E���]� �̋�U��Q�M��E���	P�M��	Q�d  ���������]� ���̋�U��j�h�h�y d�    P���SVW���1E�3�P�E�d�    �}��   �/N  ��u3��  ��  ��u�VN  3��  �M  �����L  �L��A  ��}��  �"N  3��i  ��G  ��|�=F  ��|j ��;  ����t�E  �  ��M  3��3  j�n;  ���H����H��  �} um�=H� ~X�H����H��E�    �=Է u�<  �!E  �,  �M  �E������   ��} u�=���t�  ��3��   �   �}��   �  h�   h�jh  j�/  ���E�}� tV�U�R���P�|�Q��Ѕ�t%j �U�R��  ��� �M��U��B�����j�E�P��#  ��3���3����}u
j ��  ���   �M�d�    Y_^[��]� �������������̋�U��}u��N  �EP�MQ�UR�   ��]� �������̋�U��j�h(�h�y d�    P���SVW���1E�3�P�E�d�    �e��E�   �} u�=H� u3��N  �E�    �}t�}uT�=� t�EP�MQ�UR���E�}� t�EP�MQ�UR�����E�}� u�E�    �E������E���   �EP�MQ�UR�&����E�}u=�}� u7�EPj �MQ�����URj �EP�����=� t�MQj �UR���} t�}u@�EP�MQ�UR������u�E�    �}� t�=� t�EP�MQ�UR���E��E������8�E���U��E�P�M�Q�N  ��Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]��������������̋�U���   �} t�;P  ��]�������̋�U���� � ���� ��`� ��� � �Ё �$� � �(�@� �,� � �0��� �4�� ]�����̃=�� �#s  ���\$�D$%�  =�  u�<$f�$f��f���d$��r  � �~D$f(f(�f(�fs�4f~�fT@f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�&g  ���D$��~D$f��f(�f��=�  |!=2  �fT �\�f�L$�D$����f�0fV0fT f�\$�D$���������������̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������̋T$�L$��ti3��D$��u���   r�=�� t�r  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$������̋�U��Qj j j��P�MQ�u  ���E��E���]��������̋�U��j�EP�p  ��]������������;��u���r  ̺P�1�  �P鬂  ���������z�����������������̋�U��j�hH�h�y d�    P���SVW���1E�3�P�E�d�    �Y9  �E�    �EP�9   ���E��E������   ��P9  ËE�M�d�    Y_^[��]����������̋�U������P��E����Q��E��U�;U�r�E�+E�����s3���   j�M�Q�"  ���E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M�U�;U�r"j}h�j�E�P�M�Q�Z  ���E��}� u:�U���U�E�;E�r%h�   h�j�M�Q�U�R�$  ���E��}� u3��Q�E�+E����M����U��E��E��M�Q�����UR��M���U����U��E�P�����E��]���������������̋�U��EP�"���������؃�]����̋�U��Qh�   h�jjj �  ���E��E�P�����������}� u�   ��U��    3���]���������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_��������̀�@s�� s����Ë���������������������������̋�U��E��w$������x���tRP�EQP�4   ��]ú�R�   P�E�   QP�   ��]���������������̋�U���@  ���3ŉE��ES�]VW�}S������������ǅ����    �C  ����������uS�   ���������5j j j�Wj h��  ��=   s&P������Qj�Wj h��  �օ�t�������������
ǅ�����h  �p  ����������t%���������PSQW��  �����"  2��������� ������u���  ��t�����   h  ������R������Ph  ������Q���S��  ����t-������������RWh`������P�EQ������RP���   �=j j h
  ������Qj�������Rj h��  �H�ׅ�t������j j h
  ������Pj�������Qj h��  �4�ׅ�t������������������������R�UPhVQSR����������u̋M�_^3�[�������]���������������̋�U��j�hh�h�y d�    P��$SVW���1E�3�P�E�d�    �e�3��E��E�  �M�MЍU�UԉE��M�QjPh�m@��	�   Ëe��E������E�M�d�    Y_^[��]������̋�U��j�h��h�y d�    P��$SVW���1E�3�P�E�d�    �e�3��E��E�  �M�MЋU�UԋM�M؍U�U܋M�M��E��U�RjPh�m@��	�   Ëe��E������E�M�d�    Y_^[��]����̋�U���  ���3ŉE��=����E�������E��   �8 SV��   �ȍq���A��u�+΃�-��   w{������3ɍd$ ���������A��u�Њ@��u�W������+�O�OG��u��������ȃ����Ȋ@��u�������+���O�OG��u������ȃ��_�����������SjPQ�������^[�M�3�������]����̋�U��M�h��h��d�    ]�̡d�����������̡h�����������̋�U�� � ]����̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    j角  ���E�    �E�x ��   �p��M��E�l���U��U�}� tV�E�M�;Qu�E��M�Q�P�E�P�������/�M�M��U�z uh�j jXhj��  ����u�랋M�QR�P������E�@    �E������   �j�.�  ��ËM�d�    Y_^[��]��������̋�U��} u��EP�MQ�UR�EP�MQ�*�  ]��������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�����������̋�U��j �]�̋�U���(]� ̋�U��Q���P�,�E��}� u �x�Q��E��U�R���P�0�E���]��������������̋�U���h�8�E��}� u��  3���  h �E�P� �t�h��M�Q� �x�h��U�R� �|�h��E�P� ����=t� t�=x� t�=|� t	�=�� u,�t�= �,�x��0�|��4����(����=���t�x�Q���R�0��u3���   �.  �t�P��t��x�Q��x��|�R��|����P����赌  ��u�   3��   h�A �t�Q��У���=���u	�~   3��rh  h�jh  j��
  ���E��}� t�U�R���P�|�Q��Ѕ�u	�4   3��(j �U�R�   ��� �M���U��B�����   ��]����̋�U��=���t���P���Q�����������=���t���R�4��������>�  ]������������̋�U��j�hȎh�y d�    P���SVW���1E�3�P�E�d�    h�8�E�E�@\�*�M�A    �U�B   �E�@p   �MƁ�   C�UƂK  C�E�@h�j賍  ���E�    �M�QhR�<�E������   �j�Ǎ  ���j�|�  ���E�   �E�M�Hl�U�zl u�E���Hl�U�BlP訕  ���E������   �j�p�  ��ËM�d�    Y_^[��]����������̋�U����D�E����P�����ЉE��}� u}j h�  h�jh  j�  ���E��}� tW�M�Q���R�|�P��Ѕ�t%j �M�Q�[������ �U���E��@�����j�M�Q�6  ���E�    �U�R�@�E���]�����������̋�U��Q�5����E��}� u
j�&  ���E���]�����������̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �E�E܃}� ��  �M܃y$ tj�U܋B$P�  ���M܃y, tj�U܋B,P�m  ���M܃y4 tj�U܋B4P�S  ���M܃y< tj�U܋B<P�9  ���M܃y@ tj�U܋B@P�  ���M܃yD tj�U܋BDP�  ���M܃yH tj�U܋BHP��  ���M܁y\�*tj�U܋B\P��  ��j��  ���E�    �M܋Qh�U��}� t%�E�P�H��u�}��tj�M�Q�  ���E������   �j��  ���j覊  ���E�   �U܋Bl�E�}� t4�M�Q��  ���U�;�t�}��t�E�8 u�M�Q��  ���E������   �j脊  ���j�U�R��  ���M�d�    Y_^[��]� �������������̋�U��=���tO�} u)���P�,��t���Q���R�,�ЉEj ���P�|�Q��ЋUR�����=���tj ���P�0]����������̋�U��Q�EP�MQ�UR��P�MQ�   ���E��E���]��̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�4   ���E��}� u�}� t荥  ��t
脥  �M���E���]��������̋�U��Q�EP�MQ�UR�EP�MQ�a   ���E��}� t�E��?�} u�} t	�U�   �E��%�EP荥  ����u�} t	�M�   3��뗋�]�������������̋�U��j�h�h�y d�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�9�  ���E�    �=�� vU�����9��u6�a  ��u!h|j h  hj��  ����u����    �������������E؃=Ġ�t�M�;Ġu̃=�� tu�UR�EP�M�Q�UR�EPj j�������uP�} t%�MQ�URh�j j j j ��{  ����u�� h�hlj j j j ��{  ����u��D  �U����  ��t�����u�E�   �}�v3�MQh�j j j j�{{  ����u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t h`hlj j j j�{  ����u̋M��$�MԋU�R��  ���E܃}� u�} t	�E�    �r  ���������}� tI�U��    �E��@    �M��A    �U��B�����E܋M�H�U��B   �E��@    �   ���+��;Mv���U����
����������E������;��v�������=�� t����M܉H�	�U܉���E܋����U��B    �E܋M�H�U܋E�B�M܋U�Q�E܋M�H�U܋E؉B�M܉��j�ȠR�E܃�P�������j�ȠQ�U�E܍L Q�������UR�ˠP�M܃� Q�������U܃� �U��E������   �j��  ��ËE��M�d�    Y_^[��]����̋�U��Q�} v�����3��u;Es��  �    3��K�E�E�E�MQ�UR�EP�MQ��R�EP�l������E��}� t�MQj �U�R��������E���]�������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�T������E��}� u�}� t�m�  ��t
�d�  �M���E���]��������̋�U��j�h8�h�y d�    P���SVW���1E�3�P�E�d�    j觃  ���E�    j�EP�MQ�UR�EP�MQ�B   ���E��E������   �j觃  ��ËE�M�d�    Y_^[��]��������������̋�U����E�    �E��M��} u�UR�EP�MQ�U�R�~������  �} t�}� u�EP�MQ�  ��3��  �=�� vV�����9��u6�  ��u!h|j h�  hj�{  ����u����    �������������U�=Ġ�t�E�;Ġu̃=�� ty�MQ�UR�E�P�MQ�U�R�EPj�������uR�} t%�MQ�URh�j j j j �v  ����u�� h\hlj j j j �tv  ����u�3��  �}��v`�} t)�UR�EP�M�Qhj j j j�:v  �� ��u���E�Ph�j j j j�v  ����u����  �    3��3  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URh�j j j j�u  ����u�� h`hlj j j j�u  ����u��Qj�ɠR�E�����P�  ����t1�MQhxj j j j�Zu  ����u��<�  �    3��t  �EP��  ����u!h0j h  hj�y  ����u̋U�� �U�E�xu�E�   �}� t8�M�y����u	�U�z t!h�j h#  hj�2y  ����u��d�M�Q����  ��u�E%��  ��u�E   �M���;Qs1�EPhlj j j j�nt  ����u��P�  �    3��  �} t%�U���$R�E�P�m�  ���E��}� u3��_  �#�M���$Q�U�R��  ���E��}� u3��:  3�u����������}� u|�=���s9�U𡄷+B������+��;M�v���U�����
��������E����+H������U�������;��v�������U��� �U�E��M�;Hv$�U��E�+BP�ˠQ�U��E�BP�K�����j�ȠQ�U�U�R�2������}� u�E��M�H�U��E�B�M��U�Q�E��M��H�} u/�} u�U�;U�t!hj h�  hj�9w  ����u̋M�;M�t�}� t�E���   �U��: t�E���U��B�A�8���;M�t!h�j h�  hj��v  ����u̋E��H����U��z t�E��H�U����7���;M�t!h�j h�  hj�v  ����u̋E������=�� t����E��B�	�M�����U𡔷��M��A    �U�����E��]�������̋�U��j�hX�h�y d�    P��SVW���1E�3�P�E�d�    j�}  ���E�    �EP�MQ�0   ���E������   �j�}  ��ËM�d�    Y_^[��]��̋�U��Q�=�� vU�����9��u6��  ��u!h|j h  hj�pu  ����u����    ����������} u�l  �}uOj�ɠP�M�����Q�B  ����t/�URh�"j j j j�p  ����u��w�  �    �  �=�� tDj j j �MQj �URj�������u%h�"hlj j j j �=p  ����u���  �MQ�  ����u!h0j h*  hj�wt  ����u̋E�� �E��M��Q����  ��tD�E��xt;�M��Q����  ��t*�E��xt!hX"j h0  hj�t  ����u̋�����m  j�ȠP�M���Q�  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��LPh�!j j j j�%o  ��(��u��<�U��� R�E��HQ�U��B%��  ��LQh !j j j j��n  �� ��u�j�ȠP�M��Q�E��L Q�Q  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��LPhx j j j j�kn  ��(��u��<�U��� R�E��HQ�U��B%��  ��LQh�j j j j�-n  �� ��u̋E��xue�M��y����u	�U��z t!hpj hi  hj�^r  ����u̋M��Q��$R�ʠP�M�Q��������U�R��}  ���Q  �E��xu�}u�E   �M��Q;Ut!h4j hw  hj��q  ����u̋M����+Q����������   �M��9 t�U���M��Q�P�6���;E�t!hj h�  hj�q  ����u̋U��B����M��y t�U��B�M����5���;E�t!h�j h�  hj�<q  ����u̋U������M��Q��$R�ʠP�M�Q�������U�R��|  ���(�E��@    �M��QR�ʠP�M��� Q�x�������]�̋�U��j�hx�h�y d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� u!h�j h�  hj�tp  ����u̃}� u1���  �    j h�  hh#h��o|  ������8  �=�� vV�����9��u6�u  ��u!h|j h�  hj��o  ����u����    ���������j��v  ���E�    �UR��  ����u!h0j h�  hj�o  ����u̋M�� �M��U��B%��  ��tC�M��yt:�U��B%��  ��t*�M��yt!hX"j h�  hj�@o  ����u̋E��xu�}u�E   �M��Q�U��E������   �j�Sv  ��ËE�M�d�    Y_^[��]����������̋�U��E�M���M��t�U�E��E���E;�t3���Ӹ   ]�������̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �����u
�   ��  j�cu  ���E�    ��  �E��}����   �}����   �M��MЋUЃ��UЃ}���   �E��$��\ hh%hlj j j j �i  ����u��   hD%hlj j j j �^i  ����u��dh %hlj j j j �<i  ����u��Bh�$hlj j j j �i  ����u�� h�$hlj j j j ��h  ����u��E�    ��  �E�   ����E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ��L�U���E��$j�ȠP�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qh�!j j j j �h  ��(��u��-�E�� P�M�QR�E�Ph !j j j j ��g  �� ��u��E�    j�ȠR�E�H�U�D
 P�B�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Phx j j j j �pg  ��(��u��-�U�� R�E�HQ�U�Rh�j j j j �Ag  �� ��u��E�    �M�y ��   �U�BP�ʠQ�U�� R��������ud�E�x t2�M�QR�E�HQ�U�� Rh($j j j j ��f  �� ��u��"�M�� Qh�#j j j j �f  ����u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�RhX#j j j j �]f  ��(��u��-�M�QR�E�� P�M�Qh,#j j j j �.f  �� ��u��E�    �G����E������   �j��q  ��ËE܋M�d�    Y_^[��]ÍI _Y =Y Y �X �������̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    ����E�}�t�M����  ���t	�E�    ��E�   �U܉U��}� u!h�%j hy  hj�i  ����u̃}� u0�*�  �    j hy  hh�%h�%�u  ������sj�p  ���E�    ����M�}�t7�U��t���   ��E��%��  ������    �M����E������   �j�cp  ��ËE�M�d�    Y_^[��]����������̋�U��3��} ��]Ë�U��} u3��1j j �E�� P���������u3���M�� Qj ��R�L]��������������̋�U��j�h؏h�y d�    P���SVW���1E�3�P�E�d�    3��} ���E܃}� u!h�'j h�  hj�4h  ����u̃}� u.蠋  �    j h�  hh�'h�'�/t  ���m  j� o  ���E�    �U�����E�    �	�M���M�}�}�U�E�D�    �M�U�D�    �ӡ���E���M���U��}� ��   �E��H����  |f�U��B%��  ��}V�M��Q����  �E�L����U��B%��  �U�L��E��H����  �U�D��M�A�U��J����  �U�D��W�E��x t/�M��QR�E��HQ�U�RhT'j j j j �yb  �� ��u���M�Qh0'j j j j �Xb  ����u������E����H,�U����B0�E������   �j��m  ��ËM�d�    Y_^[��]��������̋�U����E�    �E�P�M��%   �M��-  P�MQ�3  ���M���   ��]����̋�U��Q�M��E��@ �} ��   ������M��A�U��B�M��Pl��E��H�U��Ah�B�M��;�t�E��H�Qp#��u
��z  �M���U��B;�t�M��Q�Bp#��u�{  �M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ������̋�U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]���̋�U��Q�M��E���]Ë�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �E�    j��k  ���E�    h�(hlj j j j �?`  ����u̃} t�M��Uࡔ��E���M��U�}� �(  �E�;E��  �M�Q����  ��t)�E�H����  t�U�B%��  ��u�����u��  �U�z twj j�E�HQ�(�������tj�U�BP�P��t$�M�QRh�(j j j j �u_  ����u��)�M�QR�E�HQh�(j j j j �J_  ����u̋E�HQhx(j j j j �(_  ����u̋E�H����  ����   �U�BP�M�Q������  R�E�� PhD(j j j j ��^  �� ��u̃=�� t,j�U�� R�P��u�E�HQ�U�� R�������E�P�MQ��   ���   �U�zu;�E�HQ�U�� Rh(j j j j �^^  ����u̋M�Q�UR�   ���Z�E�H����  ��uI�U�BP�M�Q������  R�E�� Ph�'j j j j �^  �� ��u̋U�R�EP�\   ��������E������   �j�i  ���h�'hlj j j j �]  ����u̋M�d�    Y_^[��]���������̋�U���t���3ŉE��EP�M������E�    �	�M����M��U�z}�E�H�M���E�   �U�;U��  �EE��H �M��M��u�����t3�M��i�������   ~ �M��V���PhW  �E�P趉  ���E��hW  �M�Q�M��,���P��  ���E��}� t	�U��U���E�    �E��M��L�蛄  ��U�葄  �     �E�Ph8�M�k��1   +�R�E�k��L�Q�Ӈ  ����}*j h	  hh�(h�(j"j�=�  �R�U   �� �-�  �M��������U��D� �E�P�M�Qh�(j j j j �\  ����u̍M�� ����M�3��������]��̋�U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP�l  �E]��̋�U���8���3ŉE��E�P�u������}� u�}� u�����t7�}� t1h)hlj j j j �^[  ����u�j �N������   �3��M�3�������]����̋�U��Q����E��E���]�����������̋�U�졠�]����̋�U��Q�=� th���  ����t�EP�����/  hLh4�?  ���E��}� t�E��Gh`y ������h0h ��  ���=�� th��謌  ����tj jj ���3���]���̋�U��j j�EP�  ��]���������̋�U��jj j �  ��]�����������̋�U���vQ  �EP�R  ��h�   ����]��������������̋�U��Q����E��	�M����M��}� t�U��: tj�E��Q���������j���R����������    ����E��	�M����M��}� t�U��: tj�E��Q��������j���R���������    j���P������j���Q�p�����j���R�P�X��������    ���    �l��������P�H��u'�=��tj��Q�����������R�<��]���������������̋�U��j�h�h�y d�    P���SVW���1E�3�P�E�d�    �  �E�    �=ط�U  �Է   �E�з�} ��   ���Q��E�}� ��   ���R��E��E�    �E�EԋM؉M�   ����   �E�    �E�    �E؃��E؋M�;M�r�;����U�9u��E�;E�s�h�M؋R��E������M؉�U܋��R��EС��P��E̋M�;M�u�U�;U�t�EЉEԋMԉM�ỦU��E��E��T���h`hP�  ��hhhd�  ���=ܷ u#j��L������� t�ܷ   �����P����E������   ��} t�   Ã} t��ط   �   �MQ�V   ���M�d�    Y_^[��]�̋�U���h,)�8�E��}� th)�E�P� �E��}� t�MQ�U���]�̋�U��EP�������MQ�T]���̋�U��j��a  ��]���������������̋�U��j��a  ��]���������������̋�U��Q�u����E��E�P�I~  ���M�Q�}f  ���U�R�!Q  ���E�P�E�  ���M�Q�y�  ���U�R��  ����]������̋�U��E;Es�M�9 t�U��ЋM���M��]�������̋�U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]�̋�U���p�E�P�hh�   hD)jj@j �Y������E��}� u�����  �M�������    �	�U���@�U����   9E�s^�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B$$�M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��E����  �}� ��  �M��U��E���E��M�M��M��}�   }�U��U���E�   �E��E��E�   �	�M����M����;U���   h�   hD)jj@j �6������E��}� u����E��   �M��U���������� ����	�M���@�M��U�����   9E�sP�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��,����E�    ��E����E��M����M��U����U��E�;E���   �M��9���   �U��:���   �E����tv�U����u�M��R�d��t[�E����M���������M��U��E���
�U��E���Jh�  �U���R�`��u����`  �E��H���U��J�;����E�    �	�E����E��}��!  �M������M��U��:�t�E��8���   �M��A��}� u	�E�������U�����҃���U��E�P�\�E��}����   �}� ��   �M�Q�d�E��}� tr�U��E���M����   ��u�U��B��@�M��A��U����   ��u�E��H���U��Jh�  �E���P�`��u����R�M��Q���E��P��M��Q��@�E��P�M��������U��B�   �M��A��������R�X3���]�̋�U����E�    �	�E����E��}�@}y�M��<��� tg�U������E��	�M���@�M��U�����   9E�s�M��y t�U���R�l��j�E�����Q��������U�����    �x�����]���̋�U����=�� u�w  �E�    �L��E��}� u����e  �M����t,�E����=t	�U����U��E�P��^  ���M��T�U���juh$*jj�E���P�P������E�M����=�� u�����   �L��U��	�E�E��E��M������   �E�P�^  �����E��M����=��   j~h$*jj�E�P��������M��U�: uj���P���������    ����rj h�   h�)h�)ht)�M�Q�U�R�E�Q�![  ��P��������U���U��B���j�L�P�Z������L�    �M��    ���   3���]����̋�U����E�    �=�� u��u  �� h  h�j �ph���   ���=�� t������t����U���E���E�E�M�Q�U�Rj j �E�P�   ���}����?s�}��r����w�M��U���;E�s����dh�   hX*j�M��U���P�������E��}� u����8�M�Q�U�R�E��M���R�E�P�M�Q�6   ���U�������E����3���]���������̋�U��E�ȷ]�̋�U����E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u3҃}� �U��E���M�U����U��w�E����U�
�} t�E�M����E���E�M���U�E����E��M�Q藅  ����t/�U����M��} t�U�E���
�U���U�E����E��M��t �}� �M����U�� t�E��	�7����M��u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"uH�E�3ҹ   ���u0�}� t�U��B��"u�M����M���E�    3҃}� �U��E���E�M�U���U��t$�} t�E� \�M���M�U����M��̋U����t�}� u�M���� t�E����	u�   �}� ��   �} tQ�U��P蹃  ����t)�M�U����M���M�U����U��E����U�
�E�M����E���E�)�M��R�h�  ����t�E����E��M����E��M����E��M����M��|����} t�U� �E���E�M����E�������} t�M�    �U���U�E����U�
��]Ë�U����E�    �x�E��}� u3���   �E��E�M����t�E���E�M����u	�E���E��؋M�+M������M�j j j j �U�R�E�Pj j ��E��}� tjJh�*j�M�Q�������E�}� u�U�R�t3��Dj j �E�P�M�Q�U�R�E�Pj j ���uj�M�Q��������E�    �U�R�t�E��]��������̋�V����=��s���t�Ѓ�����r�^����������̋�V� ���=�s���t�Ѓ����r�^����������̋�U��Q�E�   j h   j �|���=� u3���   ��]���������̋�U���P����    ]���̋�U���0�E� �E�   �E���E��M����M�U��B3���EԋM�Q�U�R�  ���E�H��f�   �U�U��E�E��M��U��Q�E��H�M���U�U؃}����   �E�k��MԍT�U�E�H�MЋU��E�}� ��   �U�M��Y[  �E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=�� t h����y  ����tj�UR������M����U�[  �E��H;M�th���U�R�M����U��[  �E��M�H�U�R�E�P�e   ���U�M�I�Z  �����&�U��z�th���E�P�M����������Z  �E��M߅�t�U�R�E�P�   ���E��]��������̋�U����E�8�t%�M��E��M��U�EB3E��E��M�苶���M�Q�E��M��U�EB3E��E��M��e�����]�̋�U����E�    �E�    �=��N�@�t���%  ��t����щ���   �U�R���E��E�M�3M��M���3E�E�� 3E�E���3E�E�U�R���E�3E�E�M�3M�M�}�N�@�u	�E�O�@���U��  ��u�E�G  ��E�E�M����U��҉����]Ë�U��}csm�u�EP�MQ�   ����3�]����������̋�U���������E��}� u3���  �E��H\Q�UR��  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����v  �E��H`�M�U��E�B`�M��y�4  �P+�U��	�E����E��P+T+9M�}�U�k��E��H\�D    �ЋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]������̋�U��Q�E�E��M��;Ut�E����E��\+k�M9M�s�ڋ\+k�U9U�s
�E��;Mt3���E���]��������̋�U��j jh�+h�+h`+h   h   j �W|  ��P莼����]���������̋�U��j �EP�   ��]�����������̋�U����EP�M�������M�R�p  ����et�E���E�M�R�C}  ����u�E�Q�@  ����xu	�U���U�E��M��M���������   ��U���M���M�U��E��M�U���E��E��M��E���E��u׍M�������]Ë�U��j �EP�   ��]�����������̋�U���V�EP�M�������M���t*�E�0�M����������   ��;�t�U���U�̋E��U���U����   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M��b�������   ��;�u	�U���U�E���E�M�U����M��E����E���t�؍M������^��]���̋�U��Q�E�������Az	�E�   ��E�    �E���]�����̋�U����} t$�EP�MQ�U�R�}  ���E�M���U��P��EP�MQ�U�R�~  ���E�M���]��������������̋�U��j �EP�MQ�UR������]���̋�U���D���3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�ҁ  ��3Ƀ} ���Mă}� u!h -j h�  h�,j�D  ����u̃}� u3�g  �    j h�  h�,hx,h -�P  ���   �  3�;E��ىM�u!hX,j h�  h�,j�C  ����u̃}� u3�g  �    j h�  h�,hx,hX,�O  ���   �   �}�u�E�E���M�3҃9-�E+�3Ƀ} ��+��E��U�R�E��P�M�Q�U�3��:-��E3Ƀ} ���P��}  ���Eȃ}� t�U� �E��(�EPj �M�Q�UR�EP�MQ�UR�   ���EȋEȋM�3��8�����]����̋�U���@�E�    �E P�M��u���3Ƀ} ���M܃}� u!h -j h3  h�,j�{B  ����u̃}� u@��e  �    j h3  h�,hL.h -�vN  ���E�   �M�������E���  3�;E��ىM�u!hX,j h4  h�,j�B  ����u̃}� u@�re  �    j h4  h�,hL.hX,�N  ���E�   �M��o����E��}  3��} ����#E��	;E��ىM�u!h�-j h<  h�,j�A  ����u̃}� u@��d  � "   j h<  h�,hL.h�-�|M  ���E�"   �M�������E���  �E��t'�M3҃9-��U�U�3��} ��P�M�Q�6  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M���������   ��M����E�E�M��Ƀ���E��}�u�U�U���E�+E�M+ȉM�j h_  h�,hL.h -h-�U�R�E�P��G  ��P萵�����M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE���<���t �U����0uj�M��Q�U�R��~  ���E�    �M�������Eċ�]������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP�M��^����} }�E    3Ƀ} ���M��}� u!h -j h�  h�,j�W>  ����u̃}� u@��a  �    j h�  h�,h�.h -�RJ  ���E�   �M�������E���  3�;E��ىM�u!hX,j h�  h�,j��=  ����u̃}� u@�Na  �    j h�  h�,h�.hX,��I  ���E�   �M��K����E��g  �E�  �M��;M��ډU�u!h`.j h�  h�,j�c=  ����u̃}� u@��`  � "   j h�  h�,h�.h`.�^I  ���E�"   �M�������E���  �M��Q�4襁  %�  �� �E��U��}��  ��   �}� ��   �}�u�U�U��	�E���E�j �MQ�U�R�E��P�MQ�������E��}� t�U� �E��E��M��?����E��[  �M�Q��-u�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���Eje�MQ�  ���E��}� t!�U��Ҁ����p�E���M����M��U�� �E��E��M������E���  �M��Q�?腀  ���� ��|����U���|���U�t�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���E�M��ɀ����a�у�:�U��M��Q�4��  %�  �� ��t�����x�����t����x���u[�E� 0�M���M�U��J���� ��l�����p�����l����p���u�E�    �E�    ��EЃ��Mԃ� �EЉM���U�1�E���E�M�M��U���U�} u�E��  ��M���������   ��M����E��P���� ��d�����h�����h��� w��d��� �p  �E�   �E�    �M܋E�U���~  �E�U��E܅���   �} ~}�M��Q���� #E�#U��M���~  f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�E�U��~  �E�U��U܃�f�U܋E���E�q����M܅���   �U��R���� #E�#U��M��@~  f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���U��D�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�E���$�p�M��U���U�M��Q�4�Q}  %�  �� +E�UԉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R��{  ����0�M��U���Uj h�  �E�P�M�Q�{  �E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q�{  �Ѓ�0�E��M���Mj jd�U�R�E�P��z  �E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�T{  �ȃ�0�U�
�E���Ej j
�M�Q�U�R�oz  �E��U��E���0�M��U���U�E�  �E�    �M�������E���]��������̋�U��EP�MQ��{  ��]���������̋�U���D���3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�Rt  ��3Ƀ} ���Mă}� u!h -j h*  h�,j�6  ����u̃}� u3�Z  �    j h*  h�,h�.h -�B  ���   ��   3�;E��ىM�u!hX,j h+  h�,j�-6  ����u̃}� u3�Y  �    j h+  h�,h�.hX,�(B  ���   �   �}�u�E�E���M�3҃9-�E+E��M�Q�U��EBP�M�Q�U�3��:-��EP�p  ���Eȃ}� t�M� �E��$�URj �E�P�MQ�UR�EP�"   ���EȋEȋM�3��Ϡ����]�����������̋�U���4�E�H���M��UR�M�� ���3��} ���E�}� u!h -j h�  h�,j�5  ����u̃}� u@�rX  �    j h�  h�,h�.h -�A  ���E�   �M��o����E��  3�;U��؉E�u!hX,j h�  h�,j�4  ����u̃}� u@��W  �    j h�  h�,h�.hX,�@  ���E�   �M�������E��B  �U��t7�E3Ƀ8-��M�M��U�;Uu�E�E��E܋M��0�U܃��U܋E��  �M�M��U�:-u�E�� -�M����M��U�z j�E�P�  ���M��0�U����U���E�M�H�M��} ��   j�U�R��  ���M��r���� ���   ��E��
��U����U��E�x }]�M��t�U�B�؉E�&�M�Q��9U}�E�E���M�Q�ډŰẺE�MQ�U�R�W  ���EPj0�M�Q赝�����E�    �M������EЋ�]������������̋�U���P���3ŉE��E�    �E�E��E� �MȉM�j�U�R�E�P�MċQR�P�>p  ��3Ƀ} ���M��}� u!h -j ho  h�,j�2  ����u̃}� u3��U  �    j ho  h�,h�.h -�|>  ���   �i  3�;E��ىM�u!hX,j hp  h�,j�2  ����u̃}� u3�U  �    j hp  h�,h�.hX,�>  ���   �  �E؋H���M܋U�3��:-��E�E��}�u�M�M���U�3��:-���M+ȉM��U�R�EP�M�Q�U�R�dl  ���E��}� t�E�  �E��   �M؋Q��9U����E��M؋Q���U܃}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP�_������D�B�M���t�U���M����M���t��U��B� �EPj�M�Q�UR�EP�MQ�������M�3��<�����]��������̋�U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�
������E��{�}fu!�E P�MQ�UR�EP�MQ�c������E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ�2������E��#�U R�EP�MQ�UR�EP�MQ�������E��E���]Ë�U��j �EP�MQ�UR�EP�MQ�UR������]�������̋�U��} t#�EP�:  ����P�MQ�UUR�Eo  ��]Ë�U��Q�E�    �	�E����E��}�
s�M����R��M�����ԋ�]�̋�U���`���3ŉE��E� �E� �E� �E� �E� �E� �E���E��E���E���E���E���E���E���E���E��E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E���E���E���E���E���E���E���E���E���E���E� �E� �E� �E� �E� �E� �E� �E׀�=� t���P��E���E��M��M؋U�U��}��  4�}��  ��  �E����E��}��   ��  �M����� �$��� �E�-�  �E��}���  �M��$��� �E�   �E��/�U��]��E� �]��M��]ȍU�R�U؃���u�LQ  � "   �E�E���c  �E�   �E��/�M��]��U��]��E� �]ȍM�Q�U؃���u� Q  � !   �U�E���  �E�   �E��/�E� �]��M��]��U��]ȍE�P�U؃���u�P  � "   �M�E����  �E�   �E��/�U��]��E� �]��M��]ȍU�R�U؃���u�hP  � !   �E�E���  �E�   �E��/�M��]��U��]��E� �]ȍM�Q�U؃���u�P  � "   �U�E���3  �E�   �E��/�E� �]��M��]��U��]ȍE�P�U؃��M�E����  �E�   �E��/�U�����  �E�   �E��/�E� �]��M��]��U��]ȍE�P�U؃���u�yO  � "   �M�E���  �E�   �E��/�U��]��E� �]��M��]ȍU�R�U؃��E�E���S  �E�   �E��/�M��]��U��]��E� �]ȍM�Q�U؃���u��N  � "   �U�E���  �E�   �E��/�E� �]��M��]��U��]ȍE�P�U؃���u�N  � !   �M�E���  �E�   �E��/�U��]��E� �]��M��P�U��E� �]��M��]��U��]ȍE�P�U؃���u�8N  � !   �M�E���O  �E�   �E��/�U��]��E� �]��M��]ȍU�R�U؃���u��M  � !   �E�E���  �E�   �E��/�M��]��U��]��E� �]ȍM�Q�U؃���u�M  � !   �U�E���  �E�   �E��/�E� �]��M��]��U��]ȍE�P�U؃���u�TM  � "   �M�E���k  �E�   �E��/�U��P�E��M��]��U��]��E� �]ȍM�Q�U؃���u��L  � !   �U�E���  �E�   �E��/�E� �P�M��U��]��E� �]��M��]ȍU�R�U؃���u�L  � !   �E�E���  �E�   �E��/�M��P�U��E� �]��M��]��U��]ȍE�P�U؃���u�@L  � !   �M�E���W  �E�   �E��/�U��P�E��M��]��U��]��E� �]ȍM�Q�U؃���u��K  � !   �U�E����  �E�   �E��/�E� �P�M��U��]��E� �]��M��]ȍU�R�U؃���u�K  � !   �E�E���  �E�   �E��/�M��P�U��E� �]��M��]��U��]ȍE�P�U؃���u�,K  � !   �M�E���C  �E�   �E��/�U��]��E� �]��M��]ȍU�R�U؃���u��J  � !   �E�E����  �E�   �E�|/�M��P�U��E� �]��M��]��U��]ȍE�P�U؃���u�J  � !   �M�E���  �E�   �E��/�U��]��E� �]��M��]ȍU�R�U؃���u�8J  � !   �E�E���O  �E�   �E��/�M��]��U��]��E� �]ȍM�Q�U؃���u��I  � !   �U�E���  �E�   �E�x/�E� �M�M��U��]��E� �]��M��]ȍU�R�U؃���u�I  � !   �E�E���   �E�   �E�t/�M��M�U��E� �]��M��]��U��]ȍE�P�U؃���u�:I  � !   �M�E���T�E�   �E�p/�U��M�E��M��]��U��]��E� �]ȍM�Q�U؃���u��H  � !   �U�E���M�3�輐����]��� G� �� ߙ +� w� Κ � �� W� �� � �� [� � ��  	
�I �� �� S� �� � g� �� � [� ��  � V� ��U��j
�����3�]����������̋�U���h��  �8�P�  ���E��M���  ���  ��   ���E�$�  ���E�}� ~C�}�~�}�t�5h��  �U�R�f  ���E��   �E�P���E�$j�  ���   �M�Q�E�P���$���E�$jj��  ���}���E�$�gh  ���]��E��E������Dzh��  �U�R��  ���E��D�B�E��� th��  �M�Q��  ���E��$�"�U�R���E��$���E�$jj�[  ����]����̋�U��j
�����3�]�����������f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U��������̋�U���(  � �����������5��=�f��f��f��f��f�%�f�-ܹ����E ���E���E���������P�  �������	 ����   ��������������������H�j�aE  ��j ��h�/���=H� u
j�;E  ��h	 ���P����]��̋�U��=�� u0�EP���E�$�����$���E�$�MQj�	  ��$�!��D  � !   h��  �UR�I  ���E]�̋�S�܃������U�k�l$���   ���3ŉE��C P�KQ�SR�'  ����u)�E�����E��KQ�SR�CP�KQ�S R�E�P��  ���KQ�.
  ����|����=�� u>��|��� t5�S R���C�$�����$���C�$�CP��|���Q�  ��$�%���|���R�B	  ��h��  �C P�a  ���C�M�3�������]��[����������̋�U����E�@    �M�A    �U�B    �E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U��t�E��  ��E�H���U�J�E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U�������������M�Q���ЋE�P�M�����҃������E�H���ʋU�J�E�����Ƀ������U�B�����M�A�U�������������M�Q���ЋE�P�M��� ��҃����E�H���ʋU�J�
  �E��E���t�M�Q���E�P�M���t�U�B���M�A�U���t�E�H���U�J�E���t�M�Q���E�P�M��� t�U�B���M�A�U�%   �E�}�   w�}�   t+�}� tI�}�   t.�K�}�   t�@�M����E��1�M�������E���M�������E���M�����E��M���   �U�t5�}�   t�}�   t�1�E����U�
�"�E������U�
��E������U�
�E%�  ���M��� ��ЋE��}  tT�M�Q ���E�P �M�Q ���E�P �M�U��Y�E�H`���U�J`�E�H`���U�J`�E�M��XP�X�U�B ���M�A �U�B �����M�A �U�E� �Z�M�Q`���E�P`�M�Q`�����E�P`�M�U��YP�  �EPjj �M�Q��U�B����t�M�����E��M�Q����t�E�����U�
�E�H����t�U�����M��U�B���t�M����E��M�Q��t�E���ߋU�
�E����M�}�wb�U��$��� �E���������   �U�
�@�E���������   �U�
�(�E���������   �U�
��E��������U�
�E������M�t�}�t�}�t.�;�U�%����   �M��%�U�%����   �M���U�%�����M��}  t�U�E�@P���M�U�BP���]�� �� ݫ ū �������̋�U��j �EP�MQ�UR�EP�MQ�UR������]�������̋�U���D�E���E��M��t �U��tj��  ���E�����E��  �M��t �U��tj��  ���E�����E��s  �M���   �U���  j�  ���E%   �E��}�   w�}�   tW�}� t �}�   tv��   �}�   ��   �   �M�������z�(��]���(����]؋U�E���   �E�������z�(��]���8����]ЋM�E���Z�U�������z�8��]���(����]ȋE�E���,�M�������z�8��]���8����]��U�E���E�����E��G  �M���;  �U���/  �E�    �E��t�E�   �M���������D��   �U�R�E��� �$�  ���]�M��   �M��}�����}�E��H�]��E�   �   ���]�����Au	�E�   ��E�    �U��U��E��f�E��M��f�M��	�U����U��}����}:�E��t�}� u�E�   �M���M�U��t�E�   ��E�M���M�봃}� t�E����]�U�E����E�   �}� t
j�H  ���E�����E��M��t�U�� tj �%  ���E����E�3��}� ����]������������̋�U��� �EP��   ���E�}� t^�M�M��U�U�E�E�M�M��U�U�E �E��M$�M�h��  �U(R�{  ���E�P�[  ����u�MQ�/   ���E��"� h��  �U(R�G  ���EP�   ���E ��]�̋�U��Q�E�E��}�t�}�~ �}�~���9  � !   ��9  � "   ��]����̋�U��Q�E�    �	�E����E��}�}�M���@�;Uu�E���D����3���]���������������̋�U��Q�E�� t	�E�   �K�M��t	�E�   �:�U��t	�E�   �)�E��t	�E�   ��M��t	�E�   ��E�    �E���]�������̋�U����E�]��E�  �E��M���  �U����f�M��E���]����������̋�U��}  �u�} u�   �X�}  ��u�} u�   �B�E%�  =�  u�   �+�M���  ���  u�U����u�} t�   �3�]�����������̋�U����E��������Dz���]��E�    ��   �E%�  ��   �M����u
�} ��   �E�������]����Au	�E�   ��E�    �U�U��E��u/�M��M�U��   �t	�E���E�M��M�U����U����E%��  f�E�}� t�M�� �  f�Mj ���E�$�d������]��.j ���E�$�L������]��U���  ����-�  �E��M�U���E���]���������������̋�U��Q��}��E���]��������������̋�U��Q�}����E���]�������������̋�U�����}��E#E�M��U��#��f�E��m��E���]��̋�U����E��t
�-P��]���M��t����-P��]������U��t
�-\��]���E��t	�������؛�M�� t���]����]���������̋�U��j�h8�h�y d�    P���SVW���1E�3�P�E�d�    �e�=�� ��   �E��@tp�=h� tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe��h�    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]��������U���0���S�ٽ\�����=�� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=�� t�#  ��8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8����3  �   [�À�8�����=\� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �81�����������(1����s4�H1�,ǅr���   �01����������� 1����v�@1VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�#X  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����K   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[��������̀zuf��\���������?�f�?f��^���٭^����l1�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����l1�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����d1���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-P1��p��� ƅp���
��
�t��������̋�U��Q�E�    �p���t
j
��   ���*A  �E��}� t
j�=  ���p���tjh  @j��  ��j�D�����]Ë�U��j�W  ����tj�W  ����u#�=X�uh�   �k   ��h�   �^   ��]���������̋�U��Q�E�    �	�E����E��}�s�M��U;� :u�E���:���3���]���������������̋�U���   ���3ŉE�EP�������E��}� ��  �E�    �}�   tN�}�   tE�}t?�M�Qj j j j�  �������������� t������t���E�   ��E�   �}� ��  j��U  ����tj��U  ������   �=X���   j��\�E�}� tq�}��tk�E�    �	�U���U�}��  s%�E�M�U��J�������U�E��P��u����E� j �U�R������P�  ��P������Q�U�R����  �}�   ��  ǅ����R�������- ����  +ȉ�����������������j h  h8>h >hp=h<=h  h ���_  ��P������3�������f��  h  ������Rj ����u:j h  h8>h >h�<h�<������P������Q�}_  ��P�����������R�5_  ������<vk������P�_  ���������TA�������j h  h8>h >h<jh<������+�������������+�Q������R�Z  ��P�����j h  h8>h >h�;h�;h  h ��V  ��P��~����j h  h8>h >h ;�E�Ph  h ��`V  ��P�~����h  h�:h �� T  ���M�3��t����]���������������̋�U��E�H�]�̋�U��E�U��DV�u�     j�E�P3�NVf�
����u3�^��]ËM�U�E�QRP����t�U��MZ  f9
u֋B<��~�8PE  u��HSW�x�D$+�3�3ۅ�t�;�r	��+�;p�rC��(;�r�;�t[C�=P� u �=L� uH�  �L���t:�P���L�h�>P� 3�;�t�U�R�UVV�M�QVVVR�Ѓ� ��u	_[3�^��]ËM����u���=��1��  �M���@�U�Rh�>V�Ѕ��p  �M��R VVV�E�PWS�҅��K  �M�u���@h�U�R�Є��(  �M�;��  ��B�Ѕ���   �M���Rj �E�P�E�P�EP�E�Pj �҄���   �E;�u�E�;�wE�;�r�M���B�Ѕ�u��   �E�����   =�����   ��    Qj ��P�������   �M���RV�E�Pj j j �E�P�҄�tR+}�;>rK�M��   ;�v
;<�r@;�r��D���Mj %��� ��M��Rpj j �EP�EP�E�P�҄�t�E�   Vj ��P���M����ҋM��P@�ҋM��P8�ҋM���P(�ҋE�_[^��]��������̋�U���  ���3ŉE��=Q� t3��M�3��q����]�V�5$h�>�Q��օ���  h�?�֋���u^�M�3��mq����]�W�= h|?V�׉�������u_^�M�3��Dq����]�Shh?V�׋؅�t4h\?V�׋���t&������Pjj h ?h  ���������tV��[_3�^�M�3���p����]Í�����Q������������R������Pj h�>Qǅ����  �Ӌ�����R����V����u�������u��������u����r�Hf9�E����u�f��E����\t�\   f��E����@���+Ѓ��\����H��  �M�����>��>��E�������>�H��>�P��>�H��>�Pf��>�Hf�P������P�$[_�M�3�^��o����]�����̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�   ���E��E�    �E���]�̋�U��EP�MQ�UR�EP�MQ�UR�\  ��]���������̋�U��P  �q  ���3ŉE��E�    �E�    �} u
�   �  ƅ���� h  ������Pj �p��u8j h<  h�?h�Ch ChCh  ������Q��
  ��P�x�����������U��E�P�  ����@v]�M�Q�  ���U��D��E�j hE  h�?h�Ch(Bj�t�Q�U�������+й  +�Q�U�R�7o  ��P�>x�����} t'�EP�<  ����@v�MQ�+  ���U�DÉE��I&  ��������<&  �     �}uǅ�����A�
ǅ���� �U���t�M�������
ǅ���� �U���t�}uǅ�����A�
ǅ���� �M���tǅ�����A�
ǅ���� �} t�E�������
ǅ���� �} tǅ�����A�
ǅ���� �} t�M�������
ǅ���� �} tǅ�����A�
ǅ���� �}� t�U��������'�} t�E�������
ǅ���� �������������}� tǅ�����?�
ǅ���� �} tǅ�����A�
ǅ���� ������R������P������Q������R������P������Q������R������P������Q������R������P�M�Q�U���?Ph(Ah�  h   ������Q� (  ��D�E�}� }*j h`  h�?h�Ch�(j"j�5$  �R�M����� �%$  ��������}� }8j he  h�?h�Ch�@hd@h   ������R��  ��P�u����h  h@@������P�Yj  ��������������uj�0  ��j�V���������u�   �3��M�3��zk����]������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�   ���E��E�    �E���]�̋�U��EP�MQ�UR�EP�MQ�UR�~`  ��]���������̋�U��X"  �Am  ���3ŉE��E�    �E�    �} u
�   �  3�f������h  ������Qj ����u8j h<  h�?h�Gh Gh�<h  ������R�,T  ��P�Ct�����������E��M�Q��S  ����@v`�U�R��S  ���M��TA��U�j hE  h�?h�Gh(Bj�x�P�M�������+����  +���P�M�Q��j  ��P��s�����} t'�UR�gS  ����@v�EP�VS  ���M�TA��U���!  � ��������!  �     �}uǅ����8F�
ǅ����4F�M���t�E�������
ǅ����4F�M���t�}uǅ����F�
ǅ����4F�E���tǅ�����;�
ǅ����4F�} t�U�������
ǅ����4F�} tǅ����F�
ǅ����4F�} t�E�������
ǅ����4F�} tǅ�����E�
ǅ����4F�}� t�M��������'�} t�U�������
ǅ����4F�������������}� tǅ����<�
ǅ����4F�} tǅ�����E�
ǅ����4F������Q������R������P������Q������R������P������Q������R������P������Q������R�E�P�M���CRh8Eh�  h   ������P�[j  ��D�E�}� }*j h`  h�?h�Gh�(j"j��  �Q�؛���� �  ��������}� }8j hc  h�?h�Gh�DhHDh   ������P�Q  ��P�-q����h  h D������Q�F  ��������������uj�+,  ��j����������u�   �3��M�3��g����]�̋�U����E�    �E�    �	�E����E��}�$}Z�M��<̈́�uK�U�k���X��E��ŀ��M����M�h�  �U��Հ�P�`��u�M��̀�    3��뗸   ��]������̋�U����E�    �	�E����E��}�$}O�M��<̀� t@�U��<Մ�t3�E��ŀ��M��U�R�lj�E�P�t������M��̀�    ��E�    �	�U����U��}�$}3�E��<ŀ� t$�M��<̈́�u�U��Հ��E�M�Q�l뾋�]��̋�U��j�hX�h�y d�    P���SVW���1E�3�P�E�d�    �E�   �=� u�����j������h�   �������E�<ŀ� t
�   �   h  h�Gjj�8w�����E�}� u�'  �    3��   j
�   ���E�    �M�<̀� uDh�  �U�R�`��u"j�E�P�.�������  �    �E�    ��M�U�̀��j�E�P��������E������   �j
�e   ��ËE��M�d�    Y_^[��]������������̋�U��E�<ŀ� u�MQ��������u
j�7������U�Հ�P��]�̋�U��E�ŀ�Q��]��������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uh�Hj jh�Hj�K�������u̃}� u0�  �    j jh�HhlHh�H�I  ���   �L  �} ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U�E�Ph�   �M��Q�Pb����3҃} �U��}� uhDHj jh�Hj��������u̃}� u0��  �    j jh�HhlHhDH�  ���   �  �M�M��U�U��E��M���E���U����U��E���E��t�M����M�t�̓}� ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�La�����H��t3�t	�E�   ��E�    �M܉M�}� uh�Gj jh�Hj�k�������u̃}� u-��  � "   j jh�HhlHh�G�i  ���"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9��s
����E���M+M����U+щU؋E�Ph�   �M+M��U�D
P�e`����3���]������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+������̋�U��Q�E�    �}�wC�EP�t   ���E��}� t�*�=� u�h  �    ��MQ��  ����u����UR�  ���9  �    3���}� u�$  �    �E���]�������̋�U��Q�=� u�l���j������h�   舙�����} t�E�E���E�   �M�Qj ��R����]���������̋�U��QV�E�    �} u�4�EPj ��Q���E��}� u�DP��  �����h  �0^��]�̋�U��E���]�̋�U��Q����E��M�Q��E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR�
   ��]������̋�U��jh �j�   ��h ���P��]������̋�U���8  ���3ŉE��}�t�EP�\  ��ǅ����    jLj ������Q�]�����������U��� ����E��E�    ǅ���    ������������������������������������f������f������f������f������f������f�������������ǅ ���  �M�������U�������E�H��������U�������E�������M��������E�j ���U�R������������ u�}� u�}�t�EP�B  ���M�3��e]����]��SVW�T$�D$�L$URPQQh�� d�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�2f  �   �C�Df  �d�    ��_^[ËL$�A   �   t3�D$�H3��\��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�e  3�3�3�3�3���U��SVWj RhF� Q��6 _^[]�U�l$RQ�t$������]� �������������̋�U��Q�EP�<�M���    t�U���   P�<�M���    t�U���   P�<�M���    t�U���   P�<�M���    t�U���   P�<�E�    �	�M����M��}�m�U����E�|H��t$�M����U�|
P t�E����M�TPR�<�E����M�|L t$�U����E�|T t�M����U�D
TP�<넋M���   �´   R�<��]�̋�U��Q�} �  �EP�H�M���    t�U���   P�H�M���    t�U���   P�H�M���    t�U���   P�H�M���    t�U���   P�H�E�    �	�M����M��}�m�U����E�|H��t$�M����U�|
P t�E����M�TPR�H�E����M�|L t$�U����E�|T t�M����U�D
TP�H넋M���   �´   R�H�E��]����̋�U��Q�E���    ��   �M���   ج��   �U���    ��   �E���   �9 ��   �U���    t4�E���   �9 u&j�U���   P�w�����M���   R�i  ���E���    t4�M���   �: u&j�E���   Q�Zw�����U���   P��h  ��j�M���   R�4w����j�E���   Q� w�����U���    to�E���   �9 uaj�U���   -�   P��v����j�M���   ��   R��v����j�E���   ��   Q�v����j�U���   P�v�����M���   ��t8�U���   ���    u&�M���   R�a  ��j�E���   Q�^v�����E�    �	�U����U��}���   �E����M�|H��t:�U����E�|P t*�M����U�D
P�8 uj�M����U�D
PP��u�����M����U�|
L t�E����M�|T uA�U����E�|L u�M����U�|
T t!h�Pj h�   h`Pj���������u̋M����U�|
L t:�E����M�|T t*�U����E�LT�9 uj�U����E�LTQ�Ju���������j�UR�7u������]Ë�U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�������}� t�E�P�������}� t�M��9 u�}��t�U�R�������E��]����������̋�U��j�hx�h�y d�    P���SVW���1E�3�P�E�d�    �ie���E��E��Hp#��t	�U��zl uDj�������E�    ��P�M���lQ�������E��E������   �j���������e���Pl�U�}� u
j 裋�����E�M�d�    Y_^[��]�����������̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �d���E��E��Hp#��t�U��zl ��   j��������E�    �E��Hh�M�U�;�tI�}� t%�E�P�H��u�}��tj�M�Q�>s�����U���Bh���M�U�R�<�E������   �j��������	�E��Hh�M�}� u
j 茊�����E�M�d�    Y_^[��]����̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �E������c���E������E܋Hh�M��UR�H  ���E�E��M;H�  hN  h�Ujh   ��e�����E��}� ��  �U܋rh��   �}��E��     �M�Q�UR��  ���E؃}� ��  �E܋HhQ�H��u�U܁zh�tj�E܋HhQ��q�����U܋E��Bh�M܋QhR�<�E܋Hp���-  ������  j��������E�    �E��H���U��B���M��Q���E�    �	�E���E�}�}�M�U�E�f�TPf�M����E�    �	�E���E�}�  }�M�M�U�A������E�    �	�M���M�}�   }�U�U�E䊊  ����׋�R�H��u�=��tj��P�p�����M����U�R�<�E������   �j��������(�}��u"�}��tj�E�P�kp�����
  �    ��E�    �E؋M�d�    Y_^[��]���������������̋�U��j�h8d�    P��$���3�P�E�d�    �E�    �E�P�M������E�    � �    �}�u)� �   ���E��E������M�蝀���E��}�c�}�u)� �   ���E��E������M��n����E��N�4�}�u.� �   �M�������Q�U��E������M��8����E���E�E��E������M������EЋM�d�    Y��]������������̋�U���,���3ŉE�V�EP��������E�} u�MQ�  ��3���  �E�    �	�U����U��}��E  �E�k�0�� �;M�+  �E�    �	�U����U��}�  s�EE��@ ���E�    �	�M����M��}�s{�U�k�0�E����0��M��	�U���U�E����tN�U��B��tC�M���U��	�E����E��M��Q9U�w!�E�����UU��B��MM��A����v����U�E�B�M�A   �U�BP�  ���M�A�E�    �	�U����U��}�s�E�k�0�M��U�u�f��p$�f�DJ�ӋMQ�#  ��3��  �����} t!�}��  t�}��  t�UR����u����k  �E�P�MQ�����9  �E�    �	�U����U��}�  s�EE��@ ��M�U�Q�E�@    �}���   �MމM��	�Uԃ��UԋE����tE�U��B��t:�M���U��	�E����E��M��Q9U�w�EE��H���UU��J����E�   �	�E����E��}��   s�MM��Q���EE��P�֋M�QR�   ���M�A�U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�  ��3���= � t�EP�   ��3�����^�M�3��M����]�����������̋�U��Q�E�E��M���  �M��}�w-�U���h� �$�T� �  ��  ��  �	�  �3���]ÍI /� 6� =� D� K�  ����̋�U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �M�A    �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U�����A���E�    �	�M����M��}�   }�UU��E������  �׋�]���������̋�U���(  ���3ŉE�������P�M�QR�����-  ǅ����    ���������������������   s��������������������ƅ���� ������������������������������������tD�����������������������������������Q9�����w������Ƅ���� ���j �M�QR�E�HQ������Rh   ������Pjj �`  �� j �M�QRh   ������Ph   ������Qh   �U�BPj �]  ��$j �M�QRh   ������Ph   ������Qh   �U�BPj ��\  ��$ǅ����    ���������������������   ��   ��������U������t:�M������Q���E������P�M�������������������  �]��������M������t:�E������H�� �U������J�E�������������������  ��E�����ƀ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�U������B���M������A�������� �E�������  �X������ar?������zw6�M������Q�� �E������P�������� �U�������  ��E�����ƀ   �<����M�3���H����]����̋�U��=�� uj��K��������   3�]����������̋�U��V��   �M��UR�   �����   �0^]��������̋�U��Q�E�    �	�E����E��}�-s�M��U;��u�E�����7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]������������̋�U��Q�uV���E��}� u	�x����E�����]���������̋�U��Q�EV���E��}� u	�|����E�����]���������̋�U��E��]�̋�U��Q��P��E��}� t�MQ�U�����u3���   ��]����������̋�U��   ]����̋�U�����    ]���������������̋�U���V3��} ���E�}� uhpVj jHhVj�p�������u̃}� u-������    j jHhVh�UhpV�n�����3��   �}�v�����    3��~�} u�E   �URj ��P���E��MQ�URj��P���E��}� u:�}� @  w�M;M�w�8   ��t�U�U���DP���������&����0�E�^��]������������̋�U����E�����j j�E�Pj ��Q����t�}�u	�E�   ��E�    �E���]���������̋�U���V�E�E��} u�MQ��������   �} u�UR�������3��   �E�    �}�w)�} u�E   �EP�MQj ��R���E���EP�������:����    3��e�}� u	�=� u%�}� t��DP�������������0�E��1�MQ�c�������u�DP�`�������������03���J���^��]������̋�U��Q�E�����j j ��P�L��u�E������E���]�̋�U��Q�E�E��M�Qj �UR�EP�MQ�=]  ����]������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�y_  ����]��̋�U��E��=   vh�Vj j8h�Vj��������u̋UR�EPj �   ��]������������̋�U����EP�M��r���M����   vh�Vj jDh�Vj�)�������u̃}�|5�}�   ,�M���r��� ���   �U�Q#E�E�M��r���E��1�'�M��r������   �B�#E�E�M��sr���E���M��fr����]��̋�U���(�EP�M��lq���}�|6�}�   -�M��er������   �E�B#M�M��M��r���E��   �M��8r��P�U�����   R��a  ����t!�E��%�   �E�M�M��E� �E�   ��U�U��E� �E�   j�M���q��� �HQ�M���q����BP�M�Q�U�R�E�Pj�M��q��P��W  �� ��u�E�    �M��lq���E���M�#M�M؍M��Uq���E؋�]���������������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u��a  ��   u������r)��$��� �Ǻ   ��r����$��� �$��� ��$�t� �� 0� T� #ъ��F�G�F���G������r���$��� �I #ъ��F���G������r���$��� �#ъ���������r���$��� �I �� �� �� �� �� �� �� �� �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��� ���� �� � � �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�|� �����$�,� �I �Ǻ   ��r��+��$��� �$�|� ��� �� �� �F#шG��������r�����$�|� �I �F#шG�F���G������r�����$�|� ��F#шG�F�G�F���G�������V�������$�|� �I 0� 8� @� H� P� X� `� s� �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�|� ���� �� �� �� �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������̋�U����E�E��M����MZ  t3��;�E��M�H<�M�U�:PE  t3�� �E���E��M����  t3���   ��]�̋�U����E�MH<�M��E�    �U��B�M��T�U���E����E��M��(�M�U��B9E�s#�M�U;Qr�E�H�U�J9Ms�E���3���]�����������̋�U��j�h �h�y d�    P���SVW���1E�3�P�E�d�    �e��E�   �E�    �E�P���������u�E�    �E������E��   �M+M�M܋U�R�E�P�������E��}� u�E�    �E������E��b�M��Q$��   ���҃��U��E������E��@�E������7�E���U؋E�3�=  �����Ëe��E�    �E������E���E������M�d�    Y_^[��]��������������̋�U��h � �� �]���������̋�U��j�h �h�y d�    P���SVW���1E�3�P�E�d�    �e��K���@x�E�}� t#�E�    �U��E�������   Ëe��E������"����M�d�    Y_^[��]Ë�U��Q�5K���@|�E��}� t�U��a�����]�������������̋�U��j�h@�h�y d�    P���SVW���1E�3�P�E�d�    �e� �P��E�}� t#�E�    �U��E�������   Ëe��E�����������M�d�    Y_^[��]������������̋�U��E�$��M�(��U�,��E�0�]�������̋�U��j�h`�h�y d�    P���SVW���1E�3�P�E�d�    �E�    �E�    �E�EċMă��Mă}���   �U���d� �$�L� �E�$��MЋ�U�E؃��E��  �E�(��MЋ�U�E؃��E���   �E�,��MЋ�U�E؃��E���   �E�0��MЋ�U�E؃��E��   �H���E��}� u�����  �M��Q\R�EP�  �����EЋMЋ�U��   �x3�t	�E�   ��E�    �M��Mȃ}� u!h�Wj h�  h(Wj�<�������u̃}� u1�����    j h�  h(Wh�Wh�W�7���������4  �E�P��E�}�u3��  �}� uj�o���}� t
j ��������E�    �}t�}t�}u,�M��Q`�U܋E��@`    �}u�M��Qd�ŰE��@d�   �}u<�P+�M��	�Uԃ��UԡP+T+9E�}�M�k��U��B\�D    ���
�9C���MЉ�E������   ��}� t
j �i�����Ã}u�U��BdPj�U���
�MQ�U���}t�}t�}u�U��E܉B`�}u	�M��ỦQd3��M�d�    Y_^[��]Ë��� N� � 1� �� ��  ������̋�U��Q�E�E��M��Q;Ut�E����E��\+k�M9M�s�ً\+k�U9U�s�E��H;Mu�E���3���]����̋�U��,�P�]�������������̋�U��E�8�]�̋�U��jj �EPj �   ��]�������̋�U��j�hhd�    P�����3�P�E�d�    �EP�M��me���E�    �M�M�M��gf���P�E�L#Mu;�} t�M��If������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E؉E��E������M���e���E��M�d�    Y��]��������������̋�U����E%�����E�M#M��������   �} tj j �|W  ���U�3�t	�E�   ��E�    �M��M��}� uhhXj j1h�Wj��������u̃}� u-������    j j1h�Wh�WhhX�������   �/�} t�EP�MQ��V  ���U���EP�MQ��V  ��3���]Ë�U����EP�M���c���M���d����t/�M���d������   ~�M���d��Pj�UR�)������E��j�EP�M��d��P�]������E�M�M�M��Yd���E��]��̋�U��=p� uj�EP���������j �MQ�U�����]Ë�U���4�EP�M��,c���}   ��   �M��'d����t/�M��d������   ~�M��d��Pj�UR�l������E��j�EP�M���c��P�������Ẽ}� t,�M���c������   �E��M��M��c���E��*  ��U�U܍M��jc���E��  �M��c��� ���   ~D�M��wc��P�M�����   Q�S  ����t"�U�����   �U��E�E��E� �E�   ������� *   �M�M��E� �E�   j�M��c����BPj�M�Q�U�R�E�Ph   �M���b����QR�M���b��P�E  ��$�E�}� u�E�E؍M��b���E��A�}�u�M��MԍM��|b���E��'��U��E���ЉUЍM��]b���E���M��Pb����]������������̋�U��Q�=p� u$�}A|�}Z�E�� �E���M�M��E���j �UR���������]�����������̋�U���@���3ŉE��E�    �E�    �EP�M���`���M���a��Pj j j j �MQ�U�R�E�P��`  �� �E��MQ�U�R�Z  ���E��E���u8�}�u�E�   �M��la���E��j��}�u�E�   �M��Pa���E��N�:�M���t�E�   �M��2a���E��0��U���t�E�   �M��a���E���E�    �M�� a���E��M�3��1����]���������������̋�U���@���3ŉE��E�    �E�    �EP�M���_���M���`��Pj j j j �MQ�U�R�E�P��_  �� �E��MQ�U�R�_  ���E��E���u8�}�u�E�   �M��\`���E��j��}�u�E�   �M��@`���E��N�:�M���t�E�   �M��"`���E��0��U���t�E�   �M��`���E���E�    �M���_���E��M�3��0����]���������������̋�U����E�E��M�Q�U�3��} ���E�}� uh -j j7h@Yj���������u̃}� u0�N����    j j7h@Yh,Yh -��������   �$  3�;U��؉E�uhX,j j8h@Yj��������u̃}� u0������    j j8h@Yh,YhX,�~������   ��  �U� 3��} ����#E��;E��ىM�uh�Xj j=h@Yj��������u̃}� u0�t���� "   j j=h@Yh,Yh�X�������"   �J  3��} ���E�}� uh�Xj j>h@Yj��������u̃}� u0�����    j j>h@Yh,Yh�X�������   ��   �U��0�E����E��} ~A�M����t�E���M�U����U���E�0   �E��M��U����U��E���E빋M�� �} |>�U����5|3�M����M��U����9u�M��0�U����U���E�����U��
�E���1u�U�B���M�A�&�U��R���������P�E��P�MQ�$  ��3���]�����������̋�U���,���3ŉE��EP�M�Q�   ���U�Rj j���ċMԉ�U؉Pf�M�f�H�l  ���U�B�E�M��U��E�Pj j(hZhZh�Y�M�Q�UR�EP�Y�����P� 7�����M�U�Q�E�M�3��7-����]���̋�U����E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E��M�����U�B�E����M��U�B%   �u;�M�Q��E���   ������ыE�P�M���E�f�M�f��f�M���U��E�ЋMf�Q��]��������������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u�K  ��   u������r)��$��Ǻ   ��r����$�$�$� ��$���4`�#ъ��F�G�F���G������r���$��I #ъ��F���G������r���$��#ъ���������r���$��I ��������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��� (4H�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��	�����$�\	�I �Ǻ   ��r��+��$���$��	���	�F#шG��������r�����$��	�I �F#шG�F���G������r�����$��	��F#шG�F�G�F���G�������V�������$��	�I `	h	p	x	�	�	�	�	�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��	���	�	�	�	�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�����������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ��������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� �����̀�@s�� s����Ë�3������3�3��̀�@s�� s����Ë�3Ҁ����3�3���U��W�}3�������ك��E���8t3�����_����̋�U��j�t\����]���������������̋�U��3�]�������̋�U����E���]��E���]���������̋�U����} uht[j jdh[j蝺������u̋M�M��U�R�U�  ���E��E��H��   u$������ 	   �U��B�� �M��A����G  �-�U��B��@t"����� "   �M��Q�� �E��P����  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6�|  �� 9E�t�y|  ��@9E�u�M�Q�{  ����u�U�R��z  ���E��H��  ��   �U��E��
+Hy!h�Zj h�   h[j��������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P��l  ���E��q�}��t!�}��t�M����U���������U���E�Р�E��H�� t7jj j �U�R�?i  ���E�U�E�#E���u�M��Q�� �E��P����O�M��Q�E���E�   �M�Q�UR�E�P�2l  ���E�M�;M�t�U��B�� �M��A�����E%�   ��]����̋�U��E����U�
�E��A�]����̋�U��E����U�
�E��A��Q�]�̋�U��E����U�
�E�f�A�]���̋�S�܃������U�k�l$���   ���3ŉE��C��M��U��U�C��M��U����U��}�w@�E��$���E�   �4�E�   �+�E�   �"�E�   ��E�   ��K�   �E�    �}� ��   �U�P�K��Q�U�R�˜������ul�C�E�}�t�}�t�}�t� �M����M��U������U��C�@�]��	�M�����M��S��R�C��P�KQ�U�R�E�P��p���Q�+�����h��  �U�P�(�����ǅl���    �K�9t�=�� u�SR�Q�������l�����l��� u�C�Q负�����M�3��!����]��[ø���������U����E�    �E�E�}� |,�}�~�}�t��T��M��U�T��y�T��E��o3�t	�E�   ��E�    �U��U��}� uh�^j j9hP^j�t�������u̃}� u+������    j j9hP^h,^h�^�r����������E���]���̋�U���@���3ŉE��E�    �+���E��E�    �E�    �E�    �=@� ��   hL_�$�Eԃ}� u3��  h@_�E�P� �E��}� u3��  �M�Q��@�h0_�U�R� P��D�h_�E�P� P��H�h _�M�Q� �E��U�R��P��=P� th�^�E�P� P��L��L�;M�th�P�;U�t]�L�P��EЋP�Q��Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W�D�;M�t�D�R��Eȃ}� t�UȉE�}� t*�H�;E�t �H�Q��Eă}� t
�U�R�UĉE�@�P��E��}� t�MQ�UR�EP�M�Q�U���3��M�3������]Ë�U���4�} t�} v	�E�   ��E�    �E�E�}� uhp`j jh`j�˲������u̃}� u0�7����    j jh`h�_hp`�ɾ�����   �\  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E��M���Qh�   �U��R������3��} ���E��}� uhDHj jh`j��������u̃}� u0�n����    j jh`h�_hDH� ������   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E܋M���Qh�   �U��R��������_��t3�t	�E�   ��E�    �U؉U�}� uhh_j j h`j��������u̃}� u0�^����    j j h`h�_hh_�������   �  �M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���MԋU���Rh�   �E��P������H��t3�t	�E�   ��E�    �EЉE�}� uh�Gj j*h`j�ޯ������u̃}� u-�J���� "   j j*h`h�_h�G�ܻ�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9��s����U���E+E����M+ȉM̋U���Rh�   �E+E��M�TAR������3���]������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uhp`j jh�`j�®������u̃}� u0�.����    j jh�`h�`hp`��������   �`  �} u`3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E�M���Qh�   �U��R������3���  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P�^����3Ƀ} ���M��}� uhDHj jh�`j蔭������u̃}� u0� ����    j jh�`h�`hDH蒹�����   �2  �E�E��M�M��}�u7�U��Ef�f�
�U���M����M��U���U��t�E����E�t���}�M����t&�M;MrhHj j+h�`j��������u̋E��Mf�f��E���U����U��E���E��t�M����M�t�U���Ut���} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �E  3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E܋M���Qh�   �U��R������H��t3�t	�E�   ��E�    �U؉U�}� uh�Gj j>h�`j�ѫ������u̃}� u-�=���� "   j j>h�`h�`h�G�Ϸ�����"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9��s����M���U+U����E+EԋM���Qh�   �U+U��E�LPQ������3���]���������������̋�U��Q�E�E��M���E����E���t��E�+E������]Ë�U���(�} t�} v	�E�   ��E�    �E�E�}� uhp`j jh�Hj蛪������u̃}� u0�����    j jh�HhDahp`虶�����   �X  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E�M���Qh�   �U��R�����3��} ���E��}� uhDHj jh�Hj�ҩ������u̃}� u0�>����    j jh�HhDahDH�е�����   �  �U�U��E�E��M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P������H��t3�t	�E�   ��E�    �E܉E�}� uh�Gj jh�Hj貨������u̃}� u-����� "   j jh�HhDah�G谴�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9��s����U���E+E����M+ȉM؋U���Rh�   �E+E��M�TAR�����3���]Ë�U��} t�E�M��U���U�E]���������������̋�U��Q�} tV�E���E�M��U��}���  u�EP�������.�}���  t%3�u!h�aj h�   hXaj�w�������u̋�]����������̋�U���]��������̋�U��j�h��h�y d�    P���PP  ��  ���1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    ƅп�� h�  j ��ѿ��P�����ƅ���� h�  j ������Q�f����3�f������h�  j ������P�G����ƅЯ�� h�  j ��ѯ��Q�*�����} |�}|����*  �E�    �}��   h���<����   j h  hbh�gh`gj
h   ��п��R�EP�z  ��P�Y����h8g���} t�M�������
ǅ����(g������R��h g����п��P��h4���[���ǅ���������=  �} ��   ǅ̯��    �������ȯ�������     �UR�EPh�  h   ��Я��Q��/  ����̯����̯�� }*j h*  hbh�gh�(j"j�����R��D���� ������ȯ�����̯�� }8j h-  hbh�gh�fhd@h   ��Я��R�T�����P������}uV�} tǅ����pf�
ǅ����\fj h2  hbh�gh�e������Ph   ��п��Q�������P�����j h4  hbh�ghPe��Я��Rh   ��п��P��t  ��P������}u�M������t8j h9  hbh�gheh eh   ��п��P�t  ��P�8����j h:  hbh�gh�dh4h   ��п��Q�yt  ��P� �����} ��   ǅį��    �$���������������     ��п��P�MQ�URh�dh�  h   ������P��������į����į�� }*j hA  hbh�gh�(j"j�����Q��B���� �������������į�� }8j hD  hbh�gh�@hd@h   ������P�Y�����P� �����:j hH  hbh�ghPd��п��Qh   ������R������P������ǅ����    ǅ����    j�������Ph   ������Q������R��r  ��������j hM  hbh�gh�cj"j������P��A���� ������ t8j hO  hbh�gh�bhxbh   ������Q�%�����P�<�����=�� u�=�� �#  ǅ����    ǅ����    j�ب�����E�   �����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   �������������렃����� un�����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   ���������������E�    �   �j������Ã����� �D  �=�� t?ǅ����    ������R������P�MQ�������tǅ����   ������������������ ��   �E������t>�U�<����t1j ������P������Q�}�����P������R�E����Q���U������t������Q���U������twƅп�� �} t9j h�  hbh�gh`gj
h   ��п��Q�UR�<t  ��P��������Я��P�MQ�U��ҍ�п��#�R�MQ�UR�x������������E������   ��}uh���HË������M�d�    Y_^[�M�3��
����]�������������̋�U��j�hБh�y d�    P���\�  �  ���1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    3�f��Я��h�  j ��ү��Q�Q	����3�f������h�  j ������P�2	����ƅ���� h�  j ������Q�	����3�f��Џ��h�  j ��ҏ��P�������} |�}|����.  �E�    �}��   h���<����   j h�  hbh�mh�mj
h   ��Я��Q�UR�.�  ��P�%����h0m���} t�E������
ǅ���m�����Q��h m����Я��R��h�l���'���ǅ���������A  �} ��   ������ ��ȏ��������     �MQ�URh�  h   ��Џ��P�H�  ����̏����̏�� }*j h  hbh�mh�(j"j�����Q�<���� �w�����ȏ�����̏�� }8j h  hbh�mh`lhHDh   ��Џ��P�������P�������}uV�} tǅ���4l�
ǅ���lj h  hbh�mh`k�����Qh   ��Я��R�~�����P�����j h  hbh�mh k��Џ��Ph   ��Я��Q������P�[�����}u�U������t8j h  hbh�mh�jh�jh   ��Я��Q�������P�����j h  hbh�mh`jh�lh   ��Я��R������P�������} ��   ǅď��    ������ �����������     ��Я��Q�UR�EPhHjh   h   ������Q�-	  ����ď����ď�� }*j h  hbh�mh�(j"j茾���R�:���� �|������������ď�� }8j h  hbh�mh�DhHDh   ������R�������P�������:j h"  hbh�mh�i��Я��Ph   ������Q������P�����ǅ����    j h(  hbh�mhXij"jj�������Rh   ������Pj �{  ��P��9���� ������������ t8j h*  hbh�mh�hhThh   ������Q�`�����P�'�����=�� u�=�� �#  ǅ����    ǅ����    j�à�����E�   �����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   �렃����� un�����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   ���E�    �   �j�������Ã����� �g  �=�� t?ǅ����    ������R������P�MQ�������t������������ǅ����   ������ �  �E�������[  �U�<�����J  �E����Q�d����������t�Jj ������R������P�������P������Q�U����P����t��   �D��t��   ǅ���    j h{  hbh�mh�gj"jj�������Qh   �����R�����P�Dx  ��P�7���� ���������� t>�����Pt5j ������Q������R�+�������P������P�M����R���@����� v������������j ������Q�����R�����P�M����R���E������t������R���E������ty3�f��Я���} t9j h�  hbh�mh�mj
h   ��Я��P�MQ�}  ��P�������Џ��R�EP�M��ɍ�Я��#�Q�EP�MQ谖�����������E������   ��}uh���HË������M�d�    Y_^[�M�3��i����]�����̋�U���@���3ŉE��E�    �����E��E�    �E�    �E�    �=T� ��   hL_�$�Eԃ}� u3��  hn�E�P� �E��}� u3��  �M�Q��T�h0_�U�R� P��X�h_�E�P� P��\�h�m�M�Q� �E��U�R��d��=d� th�^�E�P� P��`��`�;M�th�d�;U�t]�`�P��EЋd�Q��Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W�X�;M�t�X�R��Eȃ}� t�UȉE�}� t*�\�;E�t �\�Q��Eă}� t
�U�R�UĉE�T�P��E��}� t�MQ�UR�EP�M�Q�U���3��M�3��D�����]Ë�U����} u3��k  3��} ���E��}� uh�nj j7hpnj蔓������u̃}� u0� ����    j j7hpnh\nh�n蒟�����   �  �} t�U;U��   �EPj �MQ�������3҃} �U��}� uhDnj j=hpnj�
�������u̃}� u-�v����    j j=hpnh\nhDn�������   �~�M;M҃��U�uhnj j>hpnj詒������u̃}� u-����� "   j j>hpnh\nhn觞�����"   ��   ��MQ�UR�EP�Ż����3���]�������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�Iu  ����]���SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ��������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� ����������̋�U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ������������XY�$����������̋�U���SVWd�5    �u��E��6j �EP�M�Q�UR��  �E�H����U�Jd�=    �]��;d�    _^[��]� ������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�4{  �� �E�_^[�E���]����̋�U����E�    �E�p7����M�3��E��U�U�E�E��M���M�d�    �E�E�d�    �UR�EP�MQ蕏  �E�E�d�    �E��]��̋�U��Q��E�H3M�����j �MQ�U�BP�M�QRj �EP�M�QR�EP�qz  �� �E��E���]����̋�U���8S�}#  u�~8�M��   ��   �E�    �Eܰ8����M�3��E��U�U�E�E�M�M�U �U��E�    �E�    �E�    �e�m�d�    �E؍E�d�    �E�   �E�E̋M�M��b	�����   �UԍE�P�M�R�Uԃ��E�    �}� td�    ��]؉d�    �	�E�d�    �E�[��]����̋�U��QS��E�H3M�����M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ�y  �� �U�z$ u�EP�MQ�6���j j j j j �U�Rh#  �~������E��]�c�k ��   [��]���̋�U��Q�} �E�HSV�pW�M�����|8����u�&����E��MN��9L���};H~���u�M���ރ} }̋E�M�UF�1�:;xw;�v�����M�_��^��[��]Ë�U��EV�u��������   �N������   ��^]����̋�U��������   ��t�M9t�@��u��   ]�3�]���̋�U��V�u���u;��   u�e���N���   ^]��T�����   �x t�H;�t���x u�^]�"����V�P^]����������U��SVWUj j h�:�u�l�  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�:d�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�:u�Q�R9Qu�   �SQ����SQ����L$�K�C�kUQPXY]Y[� �����������̋�U��} u�W  j�E�HQ������j�U�BP������j�M�QR�����j�E�HQ�����j�U�BP�����j�M�QR�}����j�E�Q�m����j�U�B P�\����j�M�Q$R�K����j�E�H(Q�:����j�U�B,P�)����j�M�Q0R�����j�E�H4Q�����j�U�BP������j�M�Q8R������j�E�H<Q������j�U�B@P������j�M�QDR�����j�E�HHQ�����j�U�BLP�����j�M�QPR�����j�E�HTQ�n����j�U�BXP�]����j�M�Q\R�L����j�E�H`Q�;����j�U�BdP�*����j�M�QhR�����j�E�HlQ�����j�U�BpP������j�M�QtR������j�E�HxQ������j�U�B|P������j�M���   R�����j�E���   Q�����j�U���   P�����j�M���   R�t����j�E���   Q�`����j�U���   P�L����j�M���   R�8����j�E���   Q�$����j�U���   P�����j�M���   R������j�E���   Q������j�U���   P������j�M���   R������j�E���   Q�����j�U���   P�����j�M���   R�����j�E���   Q�p����j�U���   P�\����j�M���   R�H����j�E���   Q�4����j�U���   P� ����j�M���   R�����j�E���   Q������j�U���   P������j�M���   R������j�E���   Q�����j�U���   P�����j�M���   R�����j�E���   Q�����j�U��   P�l����j�M��  R�X����j�E��  Q�D����j�U��  P�0����j�M��  R�����j�E��  Q�����j�U��  P������j�M��  R������j�E��   Q������j�U��$  P�����j�M��(  R�����j�E��,  Q�����j�U��0  P�|����j�M��4  R�h����j�E��8  Q�T����j�U��<  P�@����j�M��@  R�,����j�E��D  Q�����j�U��H  P�����j�M��L  R������j�E��P  Q������j�U��T  P������j�M��X  R�����j�E��\  Q�����j�U��`  P�����]�������̋�U��} u�   �E�;جtj�U�P�V�����M�Q;ܬtj�E�HQ�7�����U�B;�tj�M�QR������E�H0;�tj�U�B0P�������M�Q4;�tj�E�H4Q������]�����̋�U��} u�  �E�H;�tj�U�BP������M�Q;�tj�E�HQ������U�B;�tj�M�QR�f�����E�H;�tj�U�BP�G�����M�Q;��tj�E�HQ�(�����U�B ;��tj�M�Q R�	�����E�H$;��tj�U�B$P�������M�Q8;�tj�E�H8Q�������U�B<;�tj�M�Q<R������E�H@;�tj�U�B@P������M�QD;�tj�E�HDQ�n�����U�BH; �tj�M�QHR�O�����E�HL;$�tj�U�BLP�0����]�����������̋�U����EP�M�����M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M�����P�   ��$�E�M�����E��]���������̋�U��� �} ~,�EP�MQ�u  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$j j �UR�EP3Ƀ}( ����   Q�U$R��E��}� u3���  �}� ~63�u2�����3��u���r#h��  �M��T	R�N�����P�%������E���E�    �E�E�}� u3��  �M�Q�U�R�EP�MQj�U$R���u
�Y  �T  j j �E�P�M�Q�UR�EP���E��}� u
�,  �'  �M��   tI�}  t>�U�;U ~
�	  �  �E P�MQ�U�R�E�P�MQ�UR����u
��   ��   ��   �E��E�}� ~63�u2�����3��u��r#h��  �U�DP�G�����P�������E���E�    �M��M��}� u�|�z�U�R�E�P�M�Q�U�R�EP�MQ����u�V�T�}  u+j j j j �U�R�E�Pj �M$Q��E��}� u�'�%�#j j �U R�EP�M�Q�U�Rj �E$P��E��}� t�M�Q�������U�R�������E���]Ë�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]����������̋�U����EP�M������M$Q�U R�EP�MQ�UR�EP�MQ�M����P�"   �� �E�M��t���E��]�������������̋�U����E�    �} u�E��Q�Uj j �EP�MQ3҃}$ ��   R�EP��E�}� u3��   3�u2�}� ~,�}����w#h��  �U�DP�T�����P�+������E���E�    �M�M��}� u3��a�U���Rj �E�P�������M�Q�U�R�EP�MQj�UR��E��}� t�EP�M�Q�U�R�EP���E��M�Q��������E���]�������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh|0j jph0j�M}������u̃}� u.蹠���    j jph0h�vh|0�K���������R  �} t�} u	�E�    ��E�   �M̉MЃ}� uh�/j jsh0j��|������u̃}� u.�?����    j jsh0h�vh�/�ш���������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �,������Eă}��t�E���UU�B� �E��x }�����������]����������̋�U��� �E�����3��} ���E��}� u!h�wj h�   h0j�w{������u̃}� u1�����    j h�   h0h�wh�w�r����������  �} t�} v	�E�   ��E�    �U�U�}� u!hPwj h�   h0j��z������u̃}� u1�c����    j h�   h0h�whPw����������d  �MQ�UR�EP�MQ�URh@���������E��}� }U�E�  �}�tI�}���t@�}v:�M��9��s����U��	�E���E�M�Qh�   �U��R��������}��uu3�t	�E�   ��E�    �M�M��}� u!hwj h�   h0j��y������u̃}� u.�f���� "   j h�   h0h�whw�����������j�}� |a�}�t[�}���tR�E���;EsG�M����U+�9��s
����E���M����U+щU��E�Ph�   �M��U�D
P��������E���]���������������̋�U���,�E������E�    3��} ���E�}� u!h�wj h  h0j� y������u̃}� u1�l����    j h  h0h�wh�w�����������  �} u�} u�} u3���  �} t�} v	�E�   ��E�    �U�U��}� u!hPwj h  h0j�gx������u̃}� u1�ӛ���    j h  h0h�whPw�b���������|  �M;M��   薛����U��EP�MQ�UR�E��P�MQh@��P������E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9��s����U���E���M+ȉM�U�Rh�   �E�M�TR�%�����������8"u
�����M������  �`�ߚ����U��EP�MQ�UR�EP�MQh@��������E��UU�B� �}��u"�}�u蛚���8"u
葚���M������Y  �}� ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�H������}��uu3�t	�E�   ��E�    �E܉E�}� u!hwj hB  h0j�gv������u̃}� u.�ә��� "   j hB  h0h�whw�b�������������z�}�t\�}���tS�U���;UsH�E����M+�9��s����U���E����M+ȉM؋U�Rh�   �E��M�TR�f������}� }	�E�������E��EԋEԋ�]�������̋�U��EPj �MQ�UR�EP�MQ�@�����]�����������̋�U����EP�M��,���M��4����U���   �P�� �  �M�M������E��]������������̋�U��j �EP������]�����������̋�U��j�h��h�y d�    P��SVW���1E�3�P�E�d�    �=��tAj��{�����E�    h�h��B��������E������   �j��{����ËM�d�    Y_^[��]����������������W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋�U�����}��E�P�   ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q��  ��f�E��m���}��U�R�X   ���E�=�� tB�EP�MQ��  ���E�U�#px�E�#px;�t�E�E�   ����E�E����E��]Ë�U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]������̋�U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]��̋�U����E%�E�]��M�Q�`   ���E�U#U�E��#E�ЉU��M�;M�u�E��+�U�R�  ���E��E�P��\�����]��M�Q�   ����]�����������̋�U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]������������̋�U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]������������̋�U��h8��EP�MQ�	   ��]����̋�U���<���3ŉE�E�H
���  ���?  �M�U�B
% �  �E�M�Q�U܋E�H�M��U����E�}����u8�E�    �M�Q��  ����t	�E�    ��U�R�  ���E�   �Z  �E�P�M�Q�  ���U�U؋E�HQ�U�R�  ����t	�E���E�M�U�A+B9E�}�M�Q�*  ���E�    �E�   ��   �U�E�;Bk�M�Q�U�R�  ���E؉E�M�Q+U�UċE�P�M�Q�Z  ���U�BP�M�Q�  ���U�B��P�M�Q�1  ���E�    �E�   �~�U�E�;|B�M�Q�  ���U܁�   ��U܋E�HQ�U�R��  ���E��UJ�M��E�   �2�E�M�H�M��U܁�����U܋E�HQ�U�R�  ���E�    �E�H���    +щU��E��M���E܋M���Ɂ�   ���EԋU�z@u�E�MԉH�U�E����M�y u�U�Eԉ�E��M�3��������]��̋�U����E�    �E���E��M����M�E虃�����E�U��  �yJ���B�   +E�   �M���U��E�M��#U�t'�E�P�MQ�n   ����u�U�R�EP��   ���E�����M���E�M#��E�M���U���U��	�E���E�}�}�M�U��    ��E���]����������̋�U����E�������E��E%  �yH���@�   +ȉM����M����҉U��E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]������������̋�U����E�������E��E%  �yH���@�   +ȉM�   �M���U�E��M��R�E�P�M��U��P�V   ���E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R�   ���E��ȋE���]������̋�U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]Ë�U����E�E��M�M��E�    �	�U����U��}�}�E�M����E���E�M����M��Ӌ�]��̋�U��Q�E�    �	�E����E��}�}�M��U��    ���]���������������̋�U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]�������̋�U���V�E�������E��E%  �yH���@�E����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U��E��M���    +M�U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]��̋�U��hP��EP�MQ�i�����]����̋�U���   ���3ŉEčE��E�3�f�M��E�   �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    3҃}$ �U��}� u!h yj h�   h�xj�xe������u̃}� u0�����    j h�   h�xhtxh y�sq����3��  �M�M��U��U��	�E����E��M���� t!�E����	t�U����
t�M����u�Ƀ}�
�s  �E���M��U����U��E���x�����x����G  ��x����$��j�U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �`�M���t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�U��"�E�   � �  f�E���E�
   �M����M��  �E�   �U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �j�M���p�����p�����+��p�����p���:w8��p������j�$��j�E�   �+�E�   �"�U����U��E�   ��E�
   �E����E���  �M���1|�U���9�E�   �E����E��K�M��U$����   ��;�u	�E�   �*�E���l�����l���0t�	�E�   ��E�
   �M��M��[  �E�   ��U���E��M����M��U���0|:�E���91�}�s �Mԃ��M��U���0�E���M����M��	�U����U���E��M$����   ��
;�u	�E�   �a�U���h�����h�����+��h�����h���:w/��h�����k�$�k�E�   �"�E����E��E�   ��E�
   �M����M��w  �E�   �E�   �}� u'��U���E��M����M��U���0u�E����E�����M���U��E����E��M���0|8�U���9/�}�s'�Eԃ��E��M���0�U��
�E����E��M����M���U���d�����d�����+��d�����d���:w/��d�����dk�$�Xk�E�   �"�E����E��E�   ��E�
   �M����M��  �E�   �U���0|�E���9�E�   �M����M���E�
   �U��U��E  �E����E��M���1|�U���9�E�	   �E����E��U�M���`�����`���+t-��`���-t��`���0t�"�E�   �&�E�   �E�������E�   ��E�
   �U��U��  �E�   ��E���M��U����U��E���0u���M���1|�U���9�E�	   �E����E���E�
   �M����M��`  �U���1|�E���9�E�	   �M����M��*�U���\�����\���0t�	�E�   ��E�
   �E��E��  �E�   ǅ|���    ��M���U��E����E��M���0|:�U���91��|���k�
�M��TЉ�|�����|���P  ~ǅ|���Q  �묋�|����E���M���U��E����E��M���0|�U���9���E�
   �E����E��d�}  tN�M����M��U���X�����X���+t��X���-t��E�   �E�������E�   ��E�
   �E��E���E�
   �M����M������U�E���}� �9  �}� �/  �}� �%  �}�v+�M���|	�U����U��E�   �E����E��M����M��}� ��   �U����U��	�E����E��M����u�Eԃ��EԋM����M��ٍU�R�E�P�M�Q�3t  ���}� }�U��ډU��E�E��E��}� u	�M�M�M��}� u	�U�+U�U��}�P  ~	�E�   �B�}�����}	�E�   �0�EP�M�Q�U�R�  ��f�E�f�E�M��M�U��U�f�E�f�E��3�f�M�3�f�U��E�E؋M؉M�}� u$3�f�U�3�f�E��M�M؋U؉U�E܃��E��V�}� t(��  f�M��E�   ��E�    3�f�U�E܃��E��(�}� t"3�f�M�3�f�U��E�E؋M؉M�U܃��U܋Ef�M�f��U�E�B�M�U؉Q�E��M���Uf�B
�E܋M�3��������]Ë�Jb�b�c)def?f$g�fwg�h h�c|c�c�c  ��d�d�d  ��e�e�e  ̋�U������3ŉE��@���`�E��} u�   �} }�M�ىM�����`�U��} u3��Mf��} tr�U���T�U��E���E�M���M�}� u�׋U�k�U��U�E���� �  |#�U��E�J�M��R�U�E���E�M�M�U�R�EP�   ��눋M�3��������]�����������̋�U���L���3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��UЁ��  f�U��E��M��f�E��U���  }�E�=�  }�M�����  ~2�U���ҁ�   ��� ���E�P�M�A    �U�    �  �E�=�?  "�M�A    �U�B    �E�     ��  �M��u9f�U�f��f�U��E�H�����u�U�z u�E�8 u3ɋUf�J
�  �EЅ�uLf�M�f��f�M��U�B%���u3�M�y u*�U�: u"�E�@    �M�A    �U�    �I  �E�    �E�    �	�E����E��}���   �M���M��E�   �   +U��U��	�Eȃ��Eȃ}� ~x�MM��MċUỦU��E�L؉M��U���M���E��E�P�M�Q�U��P�"������E��}� t�M�f�T�f���E�f�T܋M����M��Ũ��U��y����E���E��<����M����?  f�M��U���~$�E�%   �u�M�Q�d  ��f�U�f��f�U����E���Qf�M�f��f�M��U���},�E؃�t	�Mԃ��MԍU�R�  ��f�E�f��f�E��̃}� t�M؃�f�M��U؁� �  �E�%�� = � u_�}��uP�E�    �}��u8�E�    �M����  u� �  f�U�f�E�f��f�E��f�M�f��f�M��	�Uރ��U��	�Eڃ��E��M����  |/�U���ҁ�   ��� ���E�P�M�A    �U�    �-�Ef�M�f��U�E܉B�M�U��Q�E��M���Uf�B
�M�3��������]����������̋�U����E���   �����ىM��U�B%   �����؉E��M���E��M�Q��U��E�P�M�Q��U��E�P��]��������������̋�U����E�H����Ɂ�   ��M��U�B�����%   ��E��M�Q��E�P�M�Q��U��E�P�M���U��E���]�����������̋�U���x���3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�E�M�M؋U�U��E�% �  f�E��M���  f�M��U���t	�E�@-��M�A �U��uM�}� uG�}� uA3��Mf��U��� �  ��҃���-�E�P�M�A�U�B0�E�@ �   �  �M���  �e  �   �Ef��}�   �u�}� tP�M؁�   @uEj j|h�zh�zh8zh,zj�U��R�[����P�u������E�@�E�    ��   �M���tW�}�   �uN�}� uHj h�   h�zh�zh�yh�yj�U��R�O[����P�������E�@�E�    �   �}�   �uK�}� uEj h�   h�zh�zh�yh�yj�M��Q��Z����P�������U�B�E�    �Cj h�   h�zh�zhHyh@yj�E��P�Z����P�z������M�A�E�    �  �U���f�U��E�%�   f�E��M���f�M��U��E����M��E�����M��E����+U��U��M���f�M�f�U�f�U��E؉E��M��M�3�f�U�j�E���P�M�Q�A������U����?  |f�E�f��f�E��M�Q�U�R��������Ef�M�f��U��tP�E�E�E�} @3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �  �}~�E   �U����?  �U�3�f�E��E�    �	�M���M�}�}�U�R�S�������}� },�E���%�   �E��	�M����M��}� ~�U�R��������E���E��M���M��	�U���U�}� ~a�E��E̋M��MЋU��UԍE�P��������M�Q��������U�R�E�P�R  ���M�Q�������U���0�E���M����M��E� 됋U����U��E���M�U����U��E��5|[�	�M����M��U��9U�r�E����9u�U��0�ًE��9E�s�M����M��Uf�f���Mf��U���M���k�	�U����U��E��9E�r�M����0u�ߋE��9E�s=3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �&�U���E�+��M�A�U�B�M�D �E܋M�3��o�����]�����������̋�U����EP�M�R�E�Q�������E��}� t0�U��Rj�E�HQ�������E��}� t�U�B���M�A�U��R�E�HQ�U�BP�M������E�}� t�M�Q���E�P�M��Q�U�BP�M�QR��������]�̋�U��j�h�h�y d�    P���SVW���1E�3�P�E�d�    �E������E������}�u!�r���     �jr��� 	   ��������  �} |�E;��s	�E�   ��E�    �MԉM܃}� uhP|j jMh�{j�N������u̃}� u<�3r���     ��q��� 	   j jMh�{h�{hP|�Z�����������C  �E���M���������D
������؉E�uh�{j jNh�{j�N������u̃}� u<�q���     �oq��� 	   j jNh�{h�{h�{�Z�����������   �UR��g  ���E�    �E���M���������D
��t �MQ�UR�EP�MQ�   ���E��U��F��p��� 	   �q���     �E������E�����3�uh{j jYh�{j�3M������u��E������   ��MQ�3h  ��ËE��U�M�d�    Y_^[��]�������̋�U����E�E��M�M��UR�e  ���E�}��u;�Bp��� 	   3�u!h{j h�   h�{j�L������u̃������   �UR�E�P�M�Q�U�R� �E��}��u#�D�E��}� t�E�P�%o�����������>�M���U���������L����U���E���������L�E��U���]��������̋�U��j�h8�h�y d�    P���SVW���1E�3�P�E�d�    �}�u�so���     �8o��� 	   ����  �} |�E;��s	�E�   ��E�    �M؉M��}� uhP|j jCh�|j�hK������u̃}� u9�o���     ��n��� 	   j jCh�|h�|hP|�[W��������/  �E���M���������D
������؉E�uh�{j jDh�|j��J������u̃}� u9�~n���     �Cn��� 	   j jDh�|h�|h�{��V��������   �UR�d  ���E�    �E���M���������D
��t�MQ�UR�EP�   ���E��?��m��� 	   ��m���     �E�����3�uh{j jOh�|j�J������u��E������   ��EP�e  ��ËE�M�d�    Y_^[��]���������������̋�U�츐<  職�����3ŉE��E�    �E�    �E�    �E��E�} u3���
  3Ƀ} ���M��}� uh�}j jmh�|j�hI������u̃}� u9�m���     ��l���    j jmh�|h|}h�}�[U��������
  �E���M���������D
$�����E��M���t	�U���uo�E��������E�uhX}j juh�|j��H������u̃}� u9�bl���     �'l���    j juh�|h|}hX}�T���������	  �U���E���������T�� tjj j �EP�_������MQ�
  ����td�U���E���������T��   tA������EԋEԋHl3҃y �U�E�P�M���U���������Q��E�}� ��  �}� t�U�����  ��E��E�    �E�    �E�EЋM�+M;M�}  �U�����  �E��3҃�
�U��E���M���������|
8 ��   �E���M���������D
4P��������u!h }j h�   h�|j�G������u̋U���E���������T4�U��EЊ�M��U���E���������D8    j�U�R�E�P�wd  �����u�  �   �M��R�y���������   �E�+E�M+ȃ�v'j�U�R�E�P�/d  �����u�O  �MЃ��M��K�U���E���������UЊ�T4�E���M���������D
8   �E����E���  �j�M�Q�U�R�c  �����u��  �EЃ��E��4�M���t	�U���u"�E�f�f�M��U�3���
���E��MЃ��M��U�����   j j j�E�Pj�M�Qj �U�R��Eȃ}� u�f  �[j �E�P�M�Q�U�R�E���M���������
P����t�M�+MM�M��U�;U�}�  ��D�E��	  �}� tl�E�   �E�j �E�P�M�Q�U�R�E���M���������
P����t!�M�;M�}�   �U���U�E����E���D�E��   �   �M���t	�U���u{�E�P��_  �����U�;�u�E����E���D�E��R�}� tG�E�   �   f�M��U�R�_  �����M�;�u�U����U��E���E���D�E���t�����  �M���U���������L��   �k  �E�    �U����?  ǅ����    ǅ����    �E������������+M;M�  ������������������������+�=�  sz������+U;Usl�����������������������������������
u!�M���M싕�����������������������������������������������q���j �M�Q������������+�R������Q�U���E���������R����t �E�E��E�������������+�9M�}���D�E��������  �E����C  �M������ǅ����    ������+U;U�  ������������������������+ʁ��  ��   ������+E;Esu������f�f����������������������������
u&�U���U�   ������f���������������������f������f����������������c���j �E�P������������+�Q������P�M���U���������Q����t �U�U��U�������������+�9E�}���D�E���������  �U������ǅ����    �E������������+M;M��  ǅt���    ������������������������+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ��x���Q������������++���P������Pj h��  ���t�����t��� u�D�E��   �   ǅp���    j �M�Q��t���+�p���R��p�����x���Q�U���E���������R����t��p���E���p�����D�E����t���;�p������t���;�p���~�������+E�E��U����Jj �M�Q�UR�EP�M���U���������Q����t�E�    �U��U��	�D�E�}� ��   �}� t0�}�u�b��� 	   �b���M���U�R��a��������V�L�E���M���������D
��@t�M���u3��%��<b���    �ab���     ������E�+E�M�3�������]Ë�U����} uht[j j.h�}j�m>������u̋t����t��U�U�j:h�}jh   輻�����E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]��������������̋�U����}�u�-a��� 	   3��   �} |�E;��s	�E�   ��E�    �M��M��}� uhP|j j(h`~j�^=������u̃}� u*��`��� 	   j j(h`~hL~hP|�\I����3���E���M���������D
��@��]���̋�U��h�]����̋�U��Q�=�� u���   ��=��}
���   h�   h�~jj���P�y���������=�� u?���   h�   h�~jj���Q�D���������=�� u
�   �   �E�    �	�U����U��}�}�E���h��M���������E�    �	�E����E��}�}f�M����U����������<�t8�M����U����������<�t�M����U����������< u�M���ǁx������3���]����̋�U����[  �з��t�fY  j���Q�H�����]���̋�U��}h�r4�}ȯw+�E-h�����P�UB�����M�Q�� �  �E�P��M�� Q��]���������������̋�U��}}#�E��P�	B�����M�Q�� �  �E�P��M�� Q��]���̋�U��}h�r4�}ȯw+�E�H������U�J�E-h�����P��A������M�� Q��]���������������̋�U��}}#�E�H������U�J�E��P�A������M�� Q��]���̋�U��Q3��} ���E��}� uh^j j)h j�:������u̃}� u+�o]���    j j)h h�~h^�F���������U�B��]���������������̋�U�졀���3�9x�����]��������������������̋�U���@�} u�} v�} t	�E�     3���  �} t	�M���������;U����E�uh�j jJhxj� 9������u̃}� u0�\���    j jJhxh`h��E�����   �\  �UR�M������M������ �x ��   �M���   ~C�} t�} v�URj �EP�:������\��� *   �\����M؍M��*����E���  �} tw3�;U��؉E�uhX,j j]hxj�I8������u̃}� u=�[��� "   j j]hxh`hX,�GD�����E�"   �M������E��x  �U�E��} t	�M�   �E�    �M������E��J  �=  �E�    �U�Rj �EP�MQj�URj �M������ �HQ��E��}� t
�}� ��   �}� ��   �D��z��   �} t�} v�URj �EP������3�t	�E�   ��E�    �U��U܃}� uhwj j{hxj�7������u̃}� u:�Z��� "   j j{hxh`hw�C�����E�"   �M������E��L�LZ��� *   �AZ����MȍM��d����E��*�} t�U�E���E�    �M��B����E���M��5�����]�̋�U��j �EP�MQ�UR�EP�������]��������������̋�U���L�E�    �} t�} u3��(  �} t�} v3��Mf�3҃} �U�}� uh��j jEh0�j��5������u̃}� u.�_Y���    j jEh0�h�h����A��������  �MQ�M��z����} �  �M��x�����z uj�E�;EsG�MM�f��Ef��MM����u�E��E؍M������E��O  �M����M��U���U뱋E��EԍM�������E��%  �  �MQ�URj��EPj	�M��������QR��E��}� t�E����EЍM������E���  �D��zt*�PX��� *   3ɋUf�
�E������M��c����E��  �E�E��M�M��	�U���U�E��M����M���tk�U����ta�M��R���P�M��R���������t@�E��H��u,��W��� *   3ҋEf��E������M�������E��#  �	�M���M��|����U�+U�U܋EP�MQ�U�R�EPj�M��������QR��E��}� u*�\W��� *   3��Mf��E������M��o����E��   �U��U��M��Y����E��   �   �M��t���� �x u�MQ��=�����E��M��%����E��j�`j j j��URj	�M��:���� �HQ��E��}� u!��V��� *   �E������M�������E�� ��U����U��M�������E���M�������]��̋�U���L�E�    �} u�} t�} t�} w	�E�    ��E�   �EĉE��}� u!h �j h�   h0�j�2������u̃}� u3�V���    j h�   h0�h�h ��>�����   ��  �} tY3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E��M���Qh�   �U��R觜�����} t	�E�     �MQ�M������U;Uv�E�E���M�M��U��U�����;E�Ƀ��M�u!h؀j h  h0�j�1������u̃}� u@�U���    j h  h0�h�h؀�=�����E�   �M������E���  �M��,���P�E�P�MQ�UR��������E�}��ux�} tX3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P�s������KT����MЍM��n����E��/  �U���U�} ��   �E�;E��   �}���   3ɋUf�
�}�tK�}���tB�}v<�E��9��s����M��	�U���U��E���Ph�   �M��Q�ך�����U�9U����E�u!h��j h  h0�j�0������u̃}� u=�xS��� "   j h  h0�h�h���<�����E�"   �M��u����E��9�U�U��E�P   3��M�Uf�DJ��} t�E�M��U��UȍM��:����Eȋ�]���̋�U��j �EP�MQ�UR�EP�MQ�`�����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uh�Hj jh`j�/������u̃}� u0�wR���    j jh`h��h�H�	;�����   �K  �} ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q������3҃} �U��}� uhDHj jh`j�F.������u̃}� u0�Q���    j jh`h��hDH�D:�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���M܋U�Rh�   �E��P��������_��t3�t	�E�   ��E�    �E؉E�}� uhh_j j h`j�;-������u̃}� u0�P���    j j h`h��hh_�99�����   �{  �U��E��
�U���M����M��U���U��t�E����E�t�̓}� ��   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���MԋU�Rh�   �E��P�������H��t3�t	�E�   ��E�    �EЉE�}� uh�Gj j*h`j�-,������u̃}� u-�O��� "   j j*h`h��h�G�+8�����"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9��s����U���E+E����M+ȉM̋U�Rh�   �E+E��M�TR�&�����3���]�������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�0   �E��j �MQ�UR�EP�MQ�   �E��E���]����������̋�U���03��} ���E�}� uh -j jfh��j��*������u̃}� u0�MN���    j jfh��h��h -��6�����   ��  3�;U��؉E�uhx�j jgh��j�*������u̃}� u0��M���    j jgh��h��hx��}6�����   �  �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���UԋE�Ph�   �M��Q莔����3҃} ��;U��؉E�uh(�j jih��j�)������u̃}� u0�*M��� "   j jih��h��h(��5�����"   ��  �}r�}$w	�E�   ��E�    �UЉU܃}� uh��j jjh��j�B)������u̃}� u0�L���    j jjh��h��h���@5�����   �O  �E�    �M�M��} t �U��-�E����E��M����M��U�ډU�E��E�E3��u�U�E3��u�E�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} v�U�;Ur��E�;Erl�M� �U�;U��؉E�u!hāj h�   h��j�8(������u̃}� u0�K��� "   j h�   h��h��hā�34�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� �������������̋�U���x���3ŉE��E�    �E�    �} t�} u3��  3��} ���EЃ}� uh��j jfh8�j�F'������u̃}� u.�J���    j jfh8�h�h���D3��������8  �UR�M�������} �.  �M������� �x ��   �M�;Msp�U�=�   ~"�EJ��� *   �E������M��`����E���  �MM��U���M��E���E��u�M��M��M��*����E��  �U����U�눋E��E��M��	����E��  �  �M��$�������   ��   �} v�UR�EP�b  ���E�M�Qj �UR�EP�MQ�URj �M������� �HQ��E��}� t3�}� u-�UU��B���u	�M����M��U��U��M��l����E���  �/I��� *   �E������M��J����E���  ��  �E�Pj �MQ�URj��EPj �M��O�����QR��E��}� t�}� u�E����E��M������E��j  �}� u�D��zt"�H��� *   �E������M�������E��7  �M�;M�  �U�Rj �M��ο��� ���   Q�U�Rj�EPj �M�豿����QR��E�}� t�}� t"�1H��� *   �E������M��L����E���  �}� |�}�v"�H��� *   �E������M������E��  �E�E�;Ev�M��M��M�������E��t  �E�    ��U����U��E����E��M�;M�}4�UU��E��LԈ
�UU����u�M��M��M�訾���E��  벋U���U������E��E��M�肾���E���   ��   �M�蝾����y ur�E�    �U�U��	�Eȃ��EȋM����t;�E�����   ~"� G��� *   �E������M������E��   �Ũ��U�벋ẺE��M�������E��t�j�M�Qj j j j��URj �M��	���� �HQ��E��}� t�}� t�F��� *   �E������M�褽���E���U����U��M�莽���E���M�聽���M�3��7�����]���̋�U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]�����̋�U���,�E�    �} t�} w�} u�} t	�E�    ��E�   �E�E��}� u!h �j h@  h8�j�"������u̃}� u3�qE���    j h@  h8�h�h �� .�����   �  �} tU�U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�������} t	�U�    �E;Ev�M�M���U�U܋E܉E�����;M�҃��U�u!h؀j hL  h8�j�!������u̃}� u3�D���    j hL  h8�h�h؀�-�����   �  �MQ�U�R�EP�MQ�������E�}��ug�} tU�U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U؋E�Ph�   �M��Q���������C��� �  �U���U�} ��   �E�;E��   �}���   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���MԋU�Rh�   �E��P�o������M9M���ډU�u!h��j hd  h8�j�������u̃}� u0�C��� "   j hd  h8�h�h���+�����"   �(�M�M��E�P   �UU��B� �} t�E�M��E���]����������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���D�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h|0j h�   h��j�������u̃}� u1�B���    j h�   h��h��h|0�*��������  �} t�} u	�E�    ��E�   �M̉MЃ}� u!h�/j h�   h��j�*������u̃}� u1�A���    j h�   h��h��h�/�%*��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �wb�����Eă}��tY�U��B���E��M��U��Q�}� |"�E��� 3ҁ��   �U��E�����U��
��E�Pj �#b�����E��}��t�E�� 3ɋU�Ef�LP��M��y }�����������]��������������̋�U���,�E������E�    3��} ���E�}� u!h�wj h9  h��j�`������u̃}� u1��?���    j h9  h��h\�h�w�[(��������&  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U��}� u!h�j h?  h��j��������u̃}� u1�3?���    j h?  h��h\�h���'��������  �M;M��   ��>����U��EP�MQ�UR�E��P�MQh ��P������E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9��s����U���E���M+ȉM�U���Rh�   �E�M�TAR�������W>���8"u
�M>���M�������  �c�9>����U��EP�MQ�UR�EP�MQh ��������E�3ҋE�Mf�TA��}��u"�}�u��=���8"u
��=���U������a  �}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P蜄�����}��ux3�t	�E�   ��E�    �U܉U�}� u!hwj hf  h��j�������u̃}� u1�'=��� "   j hf  h��h\�hw�%��������   ����|�}�t^�}���tU�M���;MsJ�U����E+�9��s����M���U����E+E؋M���Qh�   �U��E�LPQ赃�����}� }	�E�������U��UԋEԋ�]������̋�U��EPj �MQ�UR�EP�MQ�0�����]�����������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�0   �E��j �MQ�UR�EP�MQ�   �E��E���]����������̋�U���03��} ���E�}� uh -j jfh��j�1������u̃}� u0�;���    j jfh��h|�h -�/$�����   �  3�;U��؉E�uhx�j jgh��j��������u̃}� u0�;;���    j jgh��h|�hx���#�����   �  3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���EԋM���Qh�   �U��R�ځ����3��} ����;E��ىM�uh(�j jih��j�
������u̃}� u0�v:��� "   j jih��h|�h(��#�����"   ��  �}r�}$w	�E�   ��E�    �EЉE܃}� uh��j jjh��j�������u̃}� u0��9���    j jjh��h|�h���"�����   �`  �E�    �U�U��} t%�-   �M�f��U����U��E����E��M�ىM�U��U�E3��u�U�E3��u�E�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} v�M�;Mr��U�;Urn3��Mf��U�;U��؉E�u!hāj h�   h��j�{������u̃}� u0��8��� "   j h�   h��h|�hā�v!�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ��������̋�U���蓏����   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   ��   �E�H��ft4�U�z t�} uj��EP�MQ�UR��  ���   ��   �   �E�x u$�M��������!���   �E�x ��   �M�9csm�uX�U�zrO�E�x"�vC�M�Q�B�E��}� t1�M$Q�U R�EP�MQ�UR�EP�MQ�UR�U��� �E��E��0�)�E P�MQ�U$R�EP�MQ�UR�EP�MQ�   �� �   ��]�������������̋�U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U��E��E��}��|�M�U�;Q}���B���E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  蓍�����    u��  耍�����   �E�r������   �M�E�j�UR��J  ����t��<B���E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u��A���������    ty�������   �E�����ǀ�       �M�Q�UR�^  ������t�C�M�Q�  ���Ѕ�t+j�EP�4  ��h���M���  hT��M�Q�FJ  ��@���U�:csm��n  �E�x�a  �M�y �t�U�z!�t�E�x"��9  �M�y �+  �U�R�E�P�M�Q�U R�EP赃�����E���M����M��U���U�E�;E���   �M�;U��E�M�;H~�ˋU�B�E��M�Q�U���E���E�M����M��}� ��   �U�B�H���M؋U�B�H��U���E܃��E܋M؃��M؃}� ~d�U؋�EԋM�QR�E�P�M�Q��  ����u���E��U�R�E$P�M Q�U�R�E�P�M�Q�UR�EP�MQ�UR�EP�f  ��,�	���D���������M��tj�UR�  ���E�����   �M��������!���   �E�x ��   �M�QR�EP�=  ���ȅ���   蚊�����   �U�茊�����   �E��~����M���   �p����U���   �}$ u�EP�MQ��~����UR�E$P��~��j��MQ�UR�EP�  ���M�QR�s  �������M���   �����U���   �@�E�x v7�M��u*�U$R�E P�M�Q�UR�EP�MQ�UR�EP��   �� ��>��轉�����    u��>����]���������̋�U��Q�M��EP�M���G  �M�����E���]� ��������̋�U��Q�M��E�� ���M��vH  ��]��̋�U��Q�M��M�������E��t�M�Q�c�����E���]� �̋�U��Q�M��EP�M��G  �M�����E���]� ��������̋�U���V�E�8  �u�c  �҈�����    tW�Ĉ���������9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP�~~������t��   �M�y t��R=���U�R�E�P�MQ�U R�EP�������E���M����M��U����U��E�;E���   �M��U;|\�E��M;HQ�U��B�����M��Q�| t�E��H�����U��B�L�Q��u�E��H�����U��B���@t�w���j�U$R�E P�M�Qj �U��B�����M�AP�UR�EP�MQ�UR�EP��  ��,�3���^��]���������������̋�U��Q�E�x t�M�Q�B��u
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q�������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]����̋�U����E��M��U���E��}�RCC�t(�}�MOC�t�}�csm�t�@�v���ǀ�       �:���b������    ~�T����   �E�M����E�3��3���]�����̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U܋E܉E��ǅ���   �E؋M؋���E؉�E�    �M�;M��   �}��~�U�E�;B}��w:���M�Q�E�M��E�   �U�B�M�|� t%�U�E��Bh  �MQ�U�B�M�T�R�l
  �E�    ��E�P�z�����Ëe��E�    �M��M��f����E������   �)��������    ~������   �EԋUԋ���MԉËU�;Uu��9���E�M�H�M�d�    Y_^[��]Ë�U����E�E��}  t�M Q�UR�E�P�MQ�  ���}, u�UR�EP�y����MQ�U,R�y���E$�Q�UR�EP�M�Q�������U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�$   ���E��}� t�EP�M�Q�Kx����]�������̋�U��j�hВh�y d�    P���SVW���1E�3�P�E�d�    �e�E�E��E�    �M�Q��U��E�HQ�U�R�{�����E�芃�����   �E��|������   �M��n����U���   �`����M���   �E�    �E�   �E�   �U R�EP�MQ�UR�EP�ix�����E��E�    ��   �M�Q�  ��Ëe�����ǀ      �U�B�E��M�y�   �U�B%�   �ȉM��	�U�B�E��M��M��U�B�E��E�    �	�Mă��MċU�E�;BsG�M�k��U��E�;D
~3�M�k��U��E�;D
!�M�k��U��D
���E��M��U��ʉE��륋M�Q�URj �EP�������E�    �E�    �E������E�    �   �   �M�U��Q��E�P�z����������Mȉ��   ������Ủ��   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP��y������t�M�Q�UR�  ��ËEЋM�d�    Y_^[��]����������̋�U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u����ǀ     �   ��3���]���̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �e��E�    �E�x t#�M�Q�B��t�M�y u�U�%   �u3���  �M���   �t�E�E���M�Q�E�L�M��E�    �U���tXj�M�QR��=  ����t9j�E�P�=  ����t'�M��U�B��M��Q�U��P�G  ���M�����4���@  �U���txj�M�QR�k=  ����tYj�E�P�Y=  ����tG�M�QR�E�HQ�U�R�D�����E�xu"�M��9 t�U��R�E��Q��  ���U����f4���   �E�x uZj�M�QR��<  ����t>j�E�P��<  ����t,�M�QR�E��P�M�QR�g  ��P�E�P��C������ 4���[j�M�QR�<  ����tAj�E�P�~<  ����t/�M�QR�k<  ����t�E���t	�E�   ��E�   ��3���E�������   Ëe���2���E������E�M�d�    Y_^[��]Ë�U��j�h�h�y d�    P���SVW���1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ�������E��}�t�}�t+�R�U��R�E�HQ�#  ��P�U�BP�M�Q�_r���)j�U��R�E�HQ��   ��P�U�BP�M�Q�4r���E�������   Ëe���1���E������M�d�    Y_^[��]����̋�U��j�h8�h�y d�    P��SVW���1E�3�P�E�d�    �e�} t�E�8csm�t�U�M�y tL�U�B�x t@�E�    �M�Q�BP�M�QR�q���E�������E�����Ëe��1���E������M�d�    Y_^[��]�̋�U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]��������̋�U����} t��K1���} u�0���E� �E�    �	�E���E�M�U�;}m�E�H�Q���U��E�H�Q��E���M����M��U����U��}� ~4�E���M�U�BP�M�Q�U����EPR�t�������t�E���뀊E��]������������̋�U��j�h�d�    PQSVW���3�P�E�d�    �e��{�����    u��`0���E�    �$0���$�]{���M���   j j �9  �E����������E������r/���M�d�    Y_^[��]Ë�U��Q�E�    �	�E����E��M�U�;}'h��E����M�Q�L�d������t����2���]��U���SQ�E���E��EU�u�M�m��t��VW��_^��]�MU���   u�   Q�wt��]Y[�� ���̋�U���4  ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��;����E�    3Ƀ} �������������� u!h^j h  h�]j�4�������u̃����� uF�"���    j h  h�]h��h^�,����ǅ��������M�藙��������  �E�������������Q��@��   ������P�������������������t-�������t$����������������������������
ǅ����Р�������H$�����х�uV�������t-�������t$����������������������������
ǅ����Р�������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u!h�\j h  h�]j��������u̃����� uF�(!���    j h  h�]h��h�\�	����ǅ��������M��"���������  3Ƀ} �������������� u!h|0j h  h�]j�7�������u̃����� uF� ���    j h  h�]h��h|0�/	����ǅ��������M�蚗��������  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���
  ������ ��  �������� |%��������x��������8����������
ǅ����    ������������������k�	��������X�����������������   3�tǅ����   �
ǅ����    ������������������ u!h�j h`  h�]j���������u̃����� uF�4���    j h`  h�]h��h�������ǅ��������M��.���������  ��������������������  �������$�L��E�    �M�����P������R�����������   ������P�MQ������R�]  ���E��������U���U����������؉�����u!h�\j h�  h�]j���������u̃����� uF�2���    j h�  h�]h��h�\������ǅ��������M��,���������  ������R�EP������Q�  ����  �E�    �UԉU؋E؉E�M�M��E�    �E������E�    �  �������������������� ������������wK�����������$�l��E����E��,�M����M��!�U����U���E��   �E��	�M����M��  ��������*u(�EP�A�����E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�;A�����EЃ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  �����������$����E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��D
  ��������������������A������������7�  ����������$����U���0  u�E�   �E��M���  tUǅ����    �UR�?����f������������Ph   ������Q�U�R������������������ t�E�   �&�EP�?����f��|�����|����������E�   �������U��W  �EP��>������x�����x��� t��x����y u����U��E�P������E��P�M���   t&��x����B�E���x�����+����E��E�   ��E�    ��x����B�E���x�����U���  �E�%0  u�M���   �M��}��uǅ��������	�UЉ�������������p����MQ�>�����E��U���  te�}� u����E��E�   �M���l�����p�����p�������p�����t��l������t��l�������l����ɋ�l���+M����M��[�}� u	����U��E���t�����p�����p�������p�����t��t������t��t�������t����ɋ�t���+E��E��  �MQ�0=������h����r�������   3�tǅ����   �
ǅ����    ��������d�����d��� u!h8\j h�  h�]j���������u̃�d��� uF�<���    j h�  h�]h��h8\�� ����ǅ��������M��6���������  ��  �U��� t��h���f������f����h�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Bh�  h\j�UЁ�]  R�4q�����E��}� t�E��E��MЁ�]  �M���EУ   �U���U�E�H��P���X�����\����M��G���P�E�P�M�Q������R�E�P�M�Q��X���R�(�P��Ѓ��M���   t$�}� u�M������P�U�R�4�P��Ѓ���������gu*�U���   u�M��ȍ��P�E�P�0�Q��Ѓ��U����-u�M���   �M��U����U��E�P��������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�):������H�����L����   �U���   t�EP�:������H�����L����   �M��� tB�U���@t�EP�9��������H�����L�����MQ�9���������H�����L����=�U���@t�EP�r9�������H�����L�����MQ�W9����3҉�H�����L����E���@t@��L��� 7|	��H��� s,��H����ً�L����� �ډ�@�����D����E�   �E����H�����@�����L�����D����E�% �  u&�M���   u��@�����D����� ��@�����D����}� }	�E�   ��M�����M��}�   ~�E�   ��@����D���u�E�    �E��E��MЋUЃ��UЅ���@����D���t{�E��RP��D���Q��@���R��^����0��T����E��RP��D���P��@���Q�:^����@�����D�����T���9~��T����������T����E���T�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅<����M���u������R�EP��<���Qj �  ��������R�EP�M�Q�U�R�8  ���E���t$�M���u������R�EP��<���Qj0��  ���}� ��   �}� ��   ǅ$���    �U���8����E܉�4�����4�����4�������4�������   ��8���f�f������������Rj��(���P��0���Q�Ϸ������$�����8�������8�����$��� u	��0��� uǅ���������&������P�MQ��0���R��(���P�;  ���Z����������Q�UR�E�P�M�Q�  �������� |$�U���t������P�MQ��<���Rj �  ���}� tj�E�P�hw�����E�    ����������� t������tǅ����    �
ǅ����   �������� ����� ��� u!h��j h�  h�]j�4�������u̃� ��� uC����    j h�  h�]h��h���,�����ǅ��������M�藇���������������� ����M��{����� ����M�3��+X����]ÍI ������W�������.�1�<�&��I�R� �I _��0��)� ���k����������c�����~���u���l�   	
��U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�v0�����E��}��u�M�������U����M���]��������������̋�U��E�M���M��~!�UR�EP�MQ�)������U�:�u���]��������̋�U��Q�E�H��@t�U�z u�E�M�U�
�`�E�M���M��~P�U��E��MQ�UR�E�P�������M���M�U�:�u �����8*u�EP�MQj?��������렋�]����U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U������3ŉE��N@  f�E��M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M�P�U��@�E�MQ豒�����UR襒�����E�P�MQ�%������UR艒�����E��M��E�    �E�    �U�R�EP�������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U���f�U�뵋E�H�� �  u�UR�������f�E�f��f�E��؋Mf�U�f�Q
�M�3���S����]��������������̋�U��Q�} ��   �E;����   �M���U���������L����   �U���E���������<�th�=X�u<�U�U��}� t�}�t�}�t�"j j���j j���
j j���E���M�������������3�����
��� 	   ����     �����]������������̋�U����}�u��
���     �
��� 	   ����2  �} |�E;��s	�E�   ��E�    �M�M��}� u!hP|j h;  h��j���������u̃}� u<�{
���     �@
��� 	   j h;  h��h̆hP|�����������   �E���M���������D
������؉E�u!h�{j h<  h��j�S�������u̃}� u9��	���     �	��� 	   j h<  h��h̆h�{�C����������U���E�����������]��������������̋�U��j�h��h�y d�    P���SVW���1E�3�P�E�d�    �E���M��������M��E�   �U��z u_j
�������E�    �E��x u,h�  �M���Q�`��u�E�    �U��B���M��A�E������   �j
�z�����Ã}� t!�U���E���������TR���E�M�d�    Y_^[��]����������̋�U��E���M���������D
P��]��������̋�U��Q�= ��u�|  �= ��u���  �(j �E�Pj�MQ� �R����u���  �f�E��]Ë�U���$�} t�} u3���  �E���u�} t3ҋEf�3���  �MQ�M���}���M���~������   t1�M���~��� ���   th��j jGhX�j���������u̍M��~����z u*�} t�Ef��Uf�
�E�   �M��T~���E��R  �M��t~��P�E�Q�n��������   �M��T~������   ~R�M��A~��� �M;��   |=3҃} ��R�EP�M��~������   R�EPj	�M��~����QR���uB�M���}��� �M;��   r�U�B��u"�r��� *   �E������M��}���E��   �M��}������   �U�M��j}���E��k�a3��} ��P�MQj�URj	�M��u}��� �HQ���u� ��� *   �E������M��}���E���E�   �M��}���E���M���|����]������̋�U��j �EP�MQ�UR�������]���̋�U��j�hГh�y d�    P���SVW���1E�3�P�E�d�    �E�    j��������E�    �E�   �	�E����E��M�;����   �Uࡄ��<� t|�M�������H��   t"�Uࡄ���Q�  �����t	�U���U�}�|=�E�������� R�lj�E������R�k�����E������    �Y����E������   �j�a�����ËE�M�d�    Y_^[��]��������̋�U��} uj �.  ���@�EP�@   ����t����+�M�Q�� @  t�EP�}�����P��  ������3�]�������̋�U����E�    �E�E�M�Q����u|�E�H��  tn�U�E�
+H�M��}� ~Z�U�R�E�HQ�U�R������P�.�����;E�u�E�H��   t�U�B����M�A��U�B�� �M�A�E������U�E�H�
�U��B    �E���]�����̋�U��j�   ��]���������������̋�U��j�h�h�y d�    P���SVW���1E�3�P�E�d�    �E�    �E�    j�y������E�    �E�    �	�E����E��M�;����   �Uࡄ��<� ��   �M�������H��   ��   �Uࡄ���Q�U�R�������E�   �E�������B%�   te�}u%�M������P����������t	�M���M��:�} u4�Uࡄ����Q��t!�E������R���������u�E������E�    �   ��E������R�E�P�������������E������   �j������Ã}u�E����E܋M�d�    Y_^[��]���������������̋�U����  ���3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��{w���E�    3Ƀ} �������������� u!h^j h  h�]j�t�������u̃����� uF�� ���    j h  h�]h��h^�l�����ǅ@��������M���w����@�����  3��} �������������� u!h|0j h  h�]j���������u̃����� uF�U ���    j h  h�]h��h|0�������ǅ<��������M��Ow����<����r  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U���`  ������ �S  �������� |%��������x��������8�����(����
ǅ(���    ��(���������������k�	��������X�����������������   3�tǅ$���   �
ǅ$���    ��$��������������� u!h�j h`  h�]j�~�������u̃����� uF������    j h`  h�]h��h��v�����ǅ8��������M���u����8����  �������� ����� ����"  �� ����$����E�   ������Q�UR������P��  ����  �E�    �MԉM؋U؉U�E�E��E�    �E������E�    �  ������������������ ����������wL�������$��$���U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��E  ��������*u(�UR�"�����E�}� }�E����E��M��ىM���U�k�
�������LЉM���  �E�    ��  ��������*u�EP��!�����EЃ}� }�E�������M�k�
�������DЉE��  ������������������I����������.�  �������L��$�8��U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��n
  ������������������A����������7�J  ����������$�|��M���0  u	�U��� �U��E�   �EP������f�������M��� tW���������   ������ƅ���� �M��r��P�M��r��� ���   Q������R������P�?�������}�E�   �f������f�������������U��E�   �  �EP�c���������������� t�������y u����U��E�P�������E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�UЉ����������������MQ������E��U��� ��   �}� u����E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M��q��P�������Q�`������t������������������������������d�}� u	����M��E�   �U�����������������������������t���������t���������������ɋ�����+U����U��  �EP�������|����ϛ������   3�tǅ���   �
ǅ���    �������x�����x��� u!h8\j h�  h�]j�0�������u̃�x��� uF�����    j h�  h�]h��h8\�(�����ǅ4��������M��o����4����  ��  �M��� t��|���f������f����|�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Ah�  h\j�MЁ�]  Q�Q�����E��}� t�U��U��E�]  �E���EУ   �M���M�U�B��J���p�����t����M��n��P�U�R�E�P������Q�U�R�E�P��p���Q�(�R��Ѓ��E�%�   t%�}� u�M��Zn��P�M�Q�4�R��Ѓ���������gu)�M���   u�M��$n��P�U�R�0�P��Ѓ��M����-u�E�   �E��M����M��U�R�V������E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�������`�����d����   �U���   t�EP�Y������`�����d����   �M��� tB�U���@t�EP���������`�����d�����MQ�����������`�����d����=�U���@t�EP���������`�����d�����MQ�����3҉�`�����d����E���@t@��d��� 7|	��`��� s,��`����ً�d����� �ډ�X�����\����E�   �E����`�����X�����d�����\����E�% �  u&�M���   u��X�����\����� ��X�����\����}� }	�E�   ��M�����M��}�   ~�E�   ��X����\���u�E�    �������E��MЋUЃ��UЅ���X����\���t{�E��RP��\���Q��X���R�!?����0��l����E��RP��\���P��X���Q�>����X�����\�����l���9~��l����������l����E���l�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅T����M���u������R�EP��T���Qj �  ��������R�EP�M�Q�U�R��  ���E���t$�M���u������R�EP��T���Qj0�_  ���}� ��   �}� ��   �U���P����E܉�L�����L�����L�������L�����~}�M��i��P�M��i��� ���   Q��P���R������P�@�������H�����H��� ǅ���������2������Q�UR������P�Z  ����P����H�����P����j����������R�EP�M�Q�U�R��  �������� |$�E���t������Q�UR��T���Pj �Y  ���}� tj�M�Q��W�����E�    �{��������� t������tǅ���    �
ǅ���   �������D�����D��� u!h��j h�  h�]j��������u̃�D��� uC������    j h�  h�]h��h��������ǅ0��������M���g����0������������,����M���g����,����M�3��8����]� �'�Z����)�l��������������� �I ���������� �a���*�'���y����j�n� �=��3��   	
��U��E�H��@t�U�z u�E����U�
�4�EP�MQ��   ���Ё���  u�E� ������M����E�]��̋�U��E�M���M��~!�UR�EP�MQ�y������U�:�u���]��������̋�U��Q�E�H��@t�U�z u�E�M�U�
�b�E�M���M��~R�Uf�f�E��MQ�UR�E�P�������M���M�U�:�u �����8*u�EP�MQj?���������랋�]�̋�U���8���3ŉE�V�E�H��@�d  �UR腐�������t@�EP�t��������t/�MQ�c����������UR�R�������������E���E�Р�E�H$�����у�tj�EP���������t@�MQ�
��������t/�UR������������EP��������������E���E�Р�M�Q$������uh�M�Q���U��E�M��H�}� |2�U�f�Mf��U����  f�UދE����U�
f�E��  ��EP�MQ��  ���  �(  �UR�I��������t@�EP�8��������t/�MQ�'����������UR��������������E���E�Р�E��H��   ��   �URj�E�P�M�Q胒������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���UԋE�MԉH�}� |.�U��M��T��E�����   �UЋE����U�
��EP�M��T�R������EЃ}��u���  �k�|����E%��  �[�E�H���M̋U�ẺB�}� |/�M�f�Ef��M����  f�MʋU����M�f�E����UR�EP�r  ��^�M�3��d3����]ËD$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �����������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��� VW�   �Ĉ�}��E�E��M�M��} t�U���t�E� @��M�Q�U�R�E�P�M�Q�_^��]� �����̋�U��Q�M��M���   �E��t�M�Q������E���]� �̋�U��Q�M��E�� ��M��A    �U��B �E�Q�M���   �E���]� �����̋�U��Q�M��E�� ��M��A    �U��B �EP�M��   �E���]� �������̋�U��Q�M��E�;Et0�M���   �M�Q��t�E�HQ�M��m   ��U��E�H�J�E���]� �����̋�U��Q�M��E�� ��M��   ��]��̋�U����M��E��x t�M��Q�U���E����E���]���̋�U����M��} tK�EP���������E��M�Q��0�����U��B�E��x t�MQ�U�R�E��HQ��������U��B��]� �������������̋�U��Q�M��E��H��t�U��BP�0�����M��A    �U��B ��]��������̋�U��j j jj jh   @h��� �]����������̋�U��= ��t�= ��t� �P�]�����������̋�U��j�h�h�y d�    P���SVW���1E�3�P�E�d�    �E�����3��} ���E��}� uh^j j.h(�j�`�������u̃}� u+������    j j.h(�h�h^�^���������W�U�B��@t�M�A    �=�UR薈�����E�    �EP�C   ���E��E������   ��MQ������ËE�M�d�    Y_^[��]�������������̋�U����E�����3��} ���E�}� uh��j jYh(�j�z�������u̃}� u.������    j jYh(�h��h���x���������   �U�U��E��H��   ta�U�R�������E��E�P�  ���M�Q�Ո����P�  ����}	�E������$�U��z tj�E��HQ�L�����U��B    �E��@    �E���]�������̋�U��j�h8�h�y d�    P���SVW���1E�3�P�E�d�    �}�u������ 	   ����  �} |�E;��s	�E�   ��E�    �M؉M��}� uhP�j j,h��j�#�������u̃}� u.����� 	   j j,h��h��hP��!���������;  �E���M���������D
������؉E�uh��j j-h��j��������u̃}� u.����� 	   j j-h��h��h�������������   �UR�������E�    �E���M���������D
��t;�MQ�������P���u�D�E���E�    �}� u�>�����U��x���� 	   �E�����3�uh{j jEh��j���������u��E������   ��UR�������ËE�M�d�    Y_^[��]���������̋�U��� �} uht[j jdh[j�m�������u̋M�M��U�R�%������E��E��H��   u&����� 	   �U��B�� �M��A���  �c  �/�U��B��@t$����� "   �M��Q�� �E��P���  �2  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6�P����� 9E�t�C�����@9E�u�M�Q�r�������u�U�R蒀�����E��H��  �  �U��E��
+Hy!h�Zj h�   h[j��������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�r�����E��s�}��t!�}��t�M����U���������U���E�Р�E��H�� t9jj j �U�R�	o�����E��U�E�#E���u�M��Q�� �E��P���  �e�M����  �U��Bf��+�E�   �M����  f�M�U�R�E�P�M�Q��q�����E�U�;U�t�E��H�� �U��J���  ��E%��  ��]�������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_����������������̋�U��j�hX�h�y d�    P���SVW���1E�3�P�E�d�    �}�u�����     �x���� 	   ����  �} |�E;��s	�E�   ��E�    �M؉M��}� uhP|j j.h؊j証������u̃}� u9�D����     �	���� 	   j j.h؊hĊhP|����������  �E���M���������D
������؉E�uh�{j j/h؊j�"�������u̃}� u9�����     ����� 	   j j/h؊hĊh�{����������   �UR��������E�    �E���M���������D
��t�MQ�n   ���E��4����� 	   �E�����3�uh{j j9h؊j�k�������u��E������   ��MQ�k�����ËE�M�d�    Y_^[��]��̋�U��QV�EP����������t]�}u������   ��u�}u(����HD��tj��������j������;�t�UR�y�����P���t	�E�    �	�D�E��EP�`������M���U���������D �}� t�M�Q�C���������3�^��]����̋�U��} uh��j j.h8�j�@�������u̋M�Q��   tK�E�H��t@j�U�BP��C�����M�Q�������E�P�M�    �U�B    �E�@    ]��%������̍M��xT���T$�B�J�3��'%���ܐ�m)��������������̍M��HT���T$�B�J�3���$������=)��������������̋T$�B�J�3���$������)�������U����   SVW��@����0   ������(��H��hP�&����_^[���   ;������]��������U����   SVW��@����0   ������j �4����_^[���   ;��f����]��̋�U��Q3��E���]��U����   SVW��@����0   ������(����_^[���   ;������]�                                                                                                                                                                                                                                                                                                                                                                                    �� ҕ � �� � � .� D� V� h� x� �� �� �� �� �� ֖ � �� � � .� <� N� ^� �� �� �� �� ԗ � � � $� >� N� d� ~� �� ��  ޘ �� � � *� 6� H� X� f� ~� �� �� �� �� ę ֙ � � � � .� D� T� f� x� �� �� �� �� ƚ         � @        �4 Т 0� �� �         R`�                My First Plugin ize Cybernetic Genetics first plugin    cg.tiff c:\program files\maxon\cinema 4d r13\plugins\firstplugin\cgmenu.cpp �   � � � � � P  Č@ P � � � � � P                    �?~   %   res ،� %s  c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp    ��*     f:\dd\vctools\crt_bld\self_x86\crt\src\dllcrt0.c    0/               �?      �?3      3            �      0C       �       ��              fmod         �2 f� �� f� ĸ f� �� f� �� �� '� �� f� f� �� f� f:\dd\vctools\crt_bld\self_x86\crt\src\onexit.c Unknown Runtime Check Error
   Stack memory around _alloca was corrupted
 A local variable was used before it was initialized
   Stack memory was corrupted
        A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
    The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
    �xT��                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.  Run-Time Check Failure #%d - %s Unknown Module Name Unknown Filename        R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s   R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .   Stack corrupted near unknown variable   
   %.2X    Stack around _alloca corrupted  Local variable used before initialization   Stack memory corruption Cast to smaller type causing loss of data   Stack pointer corruption    ���`@        f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ e h \ t y p n a m e . c p p     p N o d e - > _ N e x t   ! =   N U L L     f:\dd\vctools\crt_bld\self_x86\crt\src\tidtable.c   FlsFree FlsSetValue FlsGetValue FlsAlloc    K E R N E L 3 2 . D L L     Client  Ignore  CRT Normal  Free    D<80(Error: memory allocation: bad memory block type.
   Invalid allocation size: %Iu bytes.
    Client hook allocation failure.
    Client hook allocation failure at file %hs line %d.
    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g h e a p . c     _ C r t C h e c k M e m o r y ( )   _ p F i r s t B l o c k   = =   p O l d B l o c k   _ p L a s t B l o c k   = =   p O l d B l o c k     f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )   Error: possible heap corruption at or near 0x%p     p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q         _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )       The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()     Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
 Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
  Client hook re-allocation failure.
 Client hook re-allocation failure at file %hs line %d.
 p U s e r D a t a   ! =   N U L L   _ p F i r s t B l o c k   = =   p H e a d   _ p L a s t B l o c k   = =   p H e a d     p H e a d - > n B l o c k U s e   = =   n B l o c k U s e   p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q         HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
   HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
       HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
 _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )     Client hook free failure.
      The Block at 0x%p was allocated by aligned routines, use _aligned_free()    _ m s i z e _ d b g     %hs located at 0x%p is %Iu bytes long.
     %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
   HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
       HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
 DAMAGED _heapchk fails with unknown return value!
  _heapchk fails with _HEAPBADPTR.
   _heapchk fails with _HEAPBADEND.
   _heapchk fails with _HEAPBADNODE.
  _heapchk fails with _HEAPBADBEGIN.
 _ C r t S e t D b g F l a g         ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )     Bad memory block found at 0x%p.
    Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
  _ C r t M e m C h e c k p o i n t   s t a t e   ! =   N U L L   Object dump complete.
  crt block at 0x%p, subtype %x, %Iu bytes long.
 normal block at 0x%p, %Iu bytes long.
  client block at 0x%p, subtype %x, %Iu bytes long.
  {%ld}   %hs(%d) :   #File Error#(%d) :  Dumping objects ->
  Data: <%s> %s
 ( * _ e r r n o ( ) )   _ p r i n t M e m B l o c k D a t a     Detected memory leaks!
 CorExitProcess  m s c o r e e . d l l   f:\dd\vctools\crt_bld\self_x86\crt\src\ioinit.c s t r c p y _ s ( * e n v ,   c c h a r s ,   p )   _ s e t e n v p         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t d e n v p . c     f:\dd\vctools\crt_bld\self_x86\crt\src\stdenvp.c    f:\dd\vctools\crt_bld\self_x86\crt\src\stdargv.c    f:\dd\vctools\crt_bld\self_x86\crt\src\a_env.c        �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �      _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )   _ s e t d e f a u l t p r e c i s i o n     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n t e l \ f p 8 . c     s i z e I n B y t e s   >   0   _ c f t o e _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c v t . c     b u f   ! =   N U L L   e+000   s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )       s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )   _ c f t o e 2 _ l   s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )     _ c f t o a _ l     _ c f t o f _ l     _ c f t o f 2 _ l   _ c f t o g _ l               �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    pow exp log10   log ��P�( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s p r i n t f . c   ( f o r m a t   ! =   N U L L )     _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh            �������             ��      �@      �               ���5�h!����?      �?  r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
         R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            �9   H9	   �8
   �8   P8   �7   �7   P7   �6   �6    6   �5   `5    5   X4    �3!    2x   �1y   �1z   �1�   �1�   |1M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y         w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )     
 
     w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )   . . .   w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )   < p r o g r a m   n a m e   u n k n o w n >     w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )     _ N M S G _ W R I T E   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 m s g . c     M S P D B 1 0 0 . D L L     r   PDBOpenValidate5    E n v i r o n m e n t D i r e c t o r y         S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 0 . 0 \ S e t u p \ V S   RegCloseKey RegQueryValueExW    RegOpenKeyExW   A D V A P I 3 2 . D L L     ... Assertion Failed    Error   Warning �?�?�?    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t . c   Microsoft Visual C++ Debug Library  _CrtDbgReport: String too long or IO Error  s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )     Debug %s!

Program: %s%s%s%s%s%s%s%s%s%s%s%s

(Press Retry to debug the application)    
Module:    
File:  
Line:  

  Expression:     

For information on how your program can cause an assertion
failure, see the Visual C++ documentation on asserts.      m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )     <program name unknown>  s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )     _ _ c r t M e s s a g e W i n d o w A   A s s e r t i o n   F a i l e d     E r r o r   W a r n i n g   �C�C�C    M i c r o s o f t   V i s u a l   C + +   D e b u g   L i b r a r y     _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r     w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )   D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n )     
 M o d u l e :     
 F i l e :     
 L i n e :     E x p r e s s i o n :           
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .     w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )   _ _ c r t M e s s a g e W i n d o w W   f:\dd\vctools\crt_bld\self_x86\crt\src\mlock.c  ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )   B u f f e r   i s   t o o   s m a l l   ( ( ( _ S r c ) ) )   ! =   N U L L     s t r c p y _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c p y _ s . i n l   ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0      Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(    �N�N�N�N�N�N�N�NxNlN`N XNPNLNHNDN@N<N8N4N(N$N NNNNNNNN\ N�M�M�M�M�MX�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�M�MpMdMPM0MM�L�L�L�LpLLL,LL�K�K�K�K�K�K�K�KtKXK8KK�J�J�JxJTJ0JJ�I�I �I�IxIXI<I    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c a l r e f . c       ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   = =   N U L L ) )     H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun f:\dd\vctools\crt_bld\self_x86\crt\src\mbctype.c    _ e x p a n d _ b a s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e x p a n d . c   p B l o c k   ! =   N U L L     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s c t y p e . c     ( u n s i g n e d ) ( c   +   1 )   < =   2 5 6     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w i n s i g . c   ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )     r a i s e   _ c o n t r o l f p _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ c o n t r l f p . c   ( " I n v a l i d   i n p u t   v a l u e " ,   0 )     p f l t   ! =   N U L L         s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )   _ f p t o s t r     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f p t o s t r . c       s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )     _ f l t o u t 2     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c f o u t . c         ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f l s b u f . c     s t r   ! =   N U L L   ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx          f:\dd\vctools\crt_bld\self_x86\crt\src\output.c     ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )     ( c h   ! =   _ T ( ' \ 0 ' ) )     (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t . c   ( s t r e a m   ! =   N U L L )     _ s e t _ e r r o r _ m o d e       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e r r m o d e . c     ( " I n v a l i d   e r r o r _ m o d e " ,   0 )   GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L         ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )   S t r i n g   i s   n o t   n u l l   t e r m i n a t e d   w c s c a t _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c a t _ s . i n l   ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0     w c s n c p y _ s   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s n c p y _ s . i n l     w c s c p y _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m a l l o c . h   ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t t . c         _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g     w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )         e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )       s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )   %s(%d) : %s     s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )   s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )         s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )     Assertion failed!   Assertion failed:       s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )   , Line  <file unknown>  Second Chance Assertion Failed: File    _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )   _ V C r t D b g R e p o r t A   w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )   _CrtDbgReport: String too long or Invalid characters in String      s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )   w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )         w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )   % s ( % d )   :   % s   w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )         w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )         w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )     A s s e r t i o n   f a i l e d !   A s s e r t i o n   f a i l e d :           w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )     
   ,   L i n e     < f i l e   u n k n o w n >     S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e         _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )   _ V C r t D b g R e p o r t W   GetUserObjectInformationA   MessageBoxA s i z e I n B y t e s   > =   c o u n t     s r c   ! =   N U L L   m e m c p y _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m c p y _ s . c   d s t   ! =   N U L L                                                                                                                                                                                                                                                                                         ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������_ v s n p r i n t f _ h e l p e r   ( " B u f f e r   t o o   s m a l l " ,   0 )       s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0   _ v s p r i n t f _ s _ l   f o r m a t   ! =   N U L L     _ v s n p r i n t f _ s _ l     	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~  _ _ s t r g t o l d 1 2 _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ i n c l u d e \ s t r g t o l d 1 2 . i n l     _ L o c a l e   ! =   N U L L   1#QNAN  s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )     1#INF   s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )   1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )     $ I 1 0 _ O U T P U T   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ x 1 0 f o u t . c     ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )   ( _ o s f i l e ( f h )   &   F O P E N )   _ l s e e k i 6 4       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k i 6 4 . c       ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )     _ w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w r i t e . c     i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )   ( ( c n t   &   1 )   = =   0 )     _ w r i t e _ n o l o c k   ( b u f   ! =   N U L L )   f:\dd\vctools\crt_bld\self_x86\crt\src\_getbuf.c    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ g e t b u f . c     _ i s a t t y       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s a t t y . c   f:\dd\vctools\crt_bld\self_x86\crt\src\_file.c  _ f i l e n o   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i l e n o . c   _ w c t o m b _ s _ l   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c t o m b . c   s i z e I n B y t e s   < =   I N T _ M A X     _ m b s t o w c s _ l _ h e l p e r     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s t o w c s . c   s   ! =   N U L L   r e t s i z e   < =   s i z e I n W o r d s     b u f f e r S i z e   < =   I N T _ M A X   _ m b s t o w c s _ s _ l   ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )   s t r c a t _ s     l e n g t h   <   s i z e I n T C h a r s   2   < =   r a d i x   & &   r a d i x   < =   3 6       s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )   s i z e I n T C h a r s   >   0     x t o a _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x t o a . c   _ w c s t o m b s _ l _ h e l p e r         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o m b s . c   p w c s   ! =   N U L L     s i z e I n B y t e s   >   r e t s i z e   _ w c s t o m b s _ s _ l   ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )   _ v s w p r i n t f _ h e l p e r   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s w p r i n t . c       s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0   _ v s n w p r i n t f _ s _ l   x t o w _ s     P�bad exception   4�p�     ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )         ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )       ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       _ o u t p u t _ s _ l   _ g e t _ o s f h a n d l e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o s f i n f o . c         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b t o w c . c   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2     _ w o u t p u t _ s _ l     ( s t r   ! =   N U L L )   csm�               �        ���� Unknown exception   C O N O U T $   f c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f c l o s e . c   _ f c l o s e _ n o l o c k     ( _ o s f i l e ( f i l e d e s )   &   F O P E N )     _ c o m m i t   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c o m m i t . c   ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )     _ c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c l o s e . c     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f r e e b u f . c   s t r e a m   ! =   N U L L         H                                                           ��Ѝ               ��           ,�<�X���    �       ����    @   ��       ����    @   t�           ��X���    8�        ����    @   ��           ����                �t�            8���            T� �           ��    T�        ����    @    �            �H�           X�d���    �       ����    @   H��        ����    @   ��           ����                ���        �y  ��  p7 �8 �: 8 h �     @*         p*     ����    ����    ����    W,     ����    ����    �����. �.     ����    ����    ����    3     ����    ����    ����9 9     ����    ����    �����9 �9     ����    ����    ����    <     ����    ����    ����    �@ ����    �@ ����    ����    ����    XC ����    �C ����    ����    ����    ,I     ����    ����    ����    �J     ����    ����    ����    1Q     ����    ����    ����    �W     ����    ����    ����    �\     ����    ����    ����    �]     ����    ����    ����    k`     ����    ����    ����    �d     ����    ����    ����    �k     ����    ����    ����Ǵ ��     ����    ����    ����    ��     ����    ����    ����    ��     ����    ����    ����    ��     ����    ����    ����    >� ����0"�   Ԑ                       ����    ����    ������ ��     ����    ����    ����Y� _�     ����    ����    ����� �     ����    ����    ����    �� ����`"�   |�                       ����    ����    ����    �'        5&����    |��    ����    �0        J.����    ����    ����    tR    ����    ����    ����    �y    ����    ����    ����    �|    P�    d�   p���    �    ����       ��    �    ����       P ����    ����    ����    ��    ��������    ����    ����    ��    ��������    ����    ������    ����    ����    ����%�+�    ����    ����    ��������@           ^�����    ����                  T�"�   d�   t�                   ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    ��        ������    ����    ����    !    ����    ����    ����    E    ����    ����    ����    ���         ښ                       �� ҕ � �� � � .� D� V� h� x� �� �� �� �� �� ֖ � �� � � .� <� N� ^� �� �� �� �� ԗ � � � $� >� N� d� ~� �� ��  ޘ �� � � *� 6� H� X� f� ~� �� �� �� �� ę ֙ � � � � .� D� T� f� x� �� �� �� �� ƚ     �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer WideCharToMultiByte  IsDebuggerPresent gMultiByteToWideChar �RaiseException  EGetProcAddress  ?LoadLibraryW  �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree GetModuleHandleW  �InterlockedIncrement  sSetLastError  GetLastError  �InterlockedDecrement  �HeapValidate  �IsBadReadPtr  ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime IsProcessorFeaturePresent �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter GetModuleFileNameW  %WriteFile �HeapFree  �HeapAlloc JGetProcessHeap  �VirtualQuery  bFreeLibrary � EnterCriticalSection  9LeaveCriticalSection  RtlUnwind hGetACP  7GetOEMCP  rGetCPInfo 
IsValidCodePage �HeapReAlloc �HeapSize  �HeapQueryInformation  �OutputDebugStringA  $WriteConsoleW �OutputDebugStringW  -LCMapStringW  iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll              1�Q    "�          � �  � �'  2�   firstplugin.dll c4d_main                                                                                                                                                                                                         �    .?AVCGMenu@@    �    .?AVCommandData@@   �    .?AVBaseData@@  Q   �    .?AVtype_info@@ u�  s�              N�@���D                                   ��������   ����   ��������    �����
                                                          ����������?         �/   �/   �/   �/   1   1!    1   �/   �/   �/   �0   �0   x/   t/    p/   �/   �/   �0   |/   �0   �0   �0   �0   �0"   �0#   �0$   �0%   �0&   �0      �      ���������              �       �D        � 0            �?<                                                                                                                                                                                                                                                                                     C       �U�U�U�U�U�U�U�U�U�U|UpUhU\UXUTUPULUHUDU@U<U8U4U0U,U$UUUUHU U�T�T�T�T�T�T�T�T�T�T�T	         �T�TxTpThT`TXTHT8T(TT T�S�S�S�S�S�S�S�S�S�S�S�S�S|SlSXSLS@S�S4S(SSS�R�R�R�R�R�R�RlR                                                                                           ��            ��            ��            ��            ��                              ج        �oxt�u���                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                     	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 0� ����        �&  �[�[����         ������������         �            .   .   Ьh�h�h�h�h�h�h�h�h�Ԭl�l�l�l�l�l�l�ج�o�q�q   ���5      @   �  �   ����             ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �    .?AVbad_exception@std@@ �    .?AVexception@std@@                .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
    ����                                                                                                                                                                                                                                                                               �                 0  �              	  H   X� Z  �      <assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel>
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPAD   T   &0�0�0+11�1�1�1�1�1�2�3{5R6W67h:o:v:}:�:�:�:�:�:�:�:�:�;L<u<�<�<h=>�>[?�?    �   #0E0�0�0;1�12�2�2�2�23*356_6�6'7�7�7�7888R8W8`8�8�8�8�8�899U9|9�9�9�9�9�9B:U:�:(;-;?;�;�;�;�;�;<<!<.<_<�<�<�<�<�<x=}=�=�=�=�=i>|>�>�>W?[?a?e?k?o?u?y??�?�?�?�?�?�?�?�?�?�?�?�?   0  ,  
0#0�0�0�0�0�01�1-2r2�2�2�2�2�293@3I3P3�3�3:4?4I4a4f4�4�4�4�4�4@6G6b6�6�627V7�7�7�7 8Q8y8�8�8�89H9M9_9�9�9�9B:|:�:�:�:�:�:;;&;8;=;O;�;�;�;�;	=='=.===D=P=W=y==�=�=�=�=�=�=�=�=�=�=�=�=�=�=�=>>>>>$>*>/>4>:>?>E>N>U>\>q>x>}>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>?&?-?P?w??�?�?�?�?�?�?�?�?�?�? @    0	00R0p0�0
11/1S1Y1`1z1�1�1�12�2+363�3�3444&4-444@4G4N4_4i4p4�4�5�5�5�5�5�566&626;6@6I6U6^66�6�6�6�67[7`7�7�788#8+848<8B8H8P8V8\8d8u8~8�8�8�89�98:=:O:/;8;A;Q;];s;;�;�;�;�;�;�;�;<<E<f<�<�<�<=%=b=n=�=�=>>�>�>�>�>�>�>�>�>�>�>�>�>?????A?]?�?�? P  (   0
0020P0Z0f0�0�0�0�0�0�0�0�0�0X1`1i1y1�1�1�1�1�1�1212=2B2r2~2�2�2�23T3Z3�3�3�344L4R4�4�4�4�45!5*5/5U5_5k5�5�5�5�5�5�5686=6O6u6�6�6�6�6�6�6�6�6�677'7M7Y7�7�7h8m88�8�8�8�89!9>9C9`9e9�9�9�9:&:/:q:�:�:;>;v;�;�;"<Q<�<�<�<�<�<�<�<�<+=7=d=i=n={=�=�=�=�=�=U>\>x>}>�>�>�>�>�>�>?[?   `  �   0'0K0V01*1B1S1�1�12;2@2i2�2�2
353W3�3�3�3�3!4}4�4�4	5�5,61666n6�677!7g7�7�7�7�7�7�7�7�7�788#8�8�8�8�8+9:9E9V9g9n9}9�9�9�9�9�9�9�9�9�9�9�9�9�9:0:=:I:Y:`:s:z:�:�:�:;;A;F;S;X;f;~;�;�;�;�;<7<^=h=�=�=�=x>�>�>�>�>�>�>�?�?�? p  �   30z0�0�0N1U1�1�1�1�1�1�1
22l2�2�2�2�2
33.33383l3{3�3�3�3�3�3�3�3�3�34U4�4�4�4A8�8�8�8�8949;9N9d9k9~9�9�9�9�9�9�9:�:�:�:;m;(<3<@<H<W<l<x<�<�<�<�<�=�=�=A?T?�?�?�?   �  d   �2�2�2333<3H3u3z33n4z4�4�4�4�4�45!5&5h5t5�5�5�5�6�6�6�6�7�8�8�8�8�899@9E9J9�9�9�9�9�9 �  �   	0T0`0�0�0�0�0�0�0�0�0�1�12!2&2X2d2�2�2�24h4t4�4�4�4�4�4	555�7�7�7�7t8|8�8�8�8�8�89Q9�9�95:�:�:�:$;a;�;�;<e<�<�<I=T=�=�=>>]>h>�>�>? ?q?�?�? �  �   0e0�0
1`1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�394>45"5(5.545:5A5H5O5V5]5d5k5s5{5�5�5�5�5�5�5�5�5�5�5�5�5�5�566'6�6�6#;�;�<�<�<�<�=�=�=�=> >C>N>�> �  �   �0144,4h4m44�4�4�4T5�56�6�6�6�6�6�6�7P8�8l9�9�9:g:s:�:I;X;�;�;�; <%<*</<9<m<}<�<�<�<�<�<�<�<9=>=C=H=R=o=t=y=�=�=�=�=>$>�>�>�>�>�>�>�>?�?�?   �  $  \0c0�0�0�0�0�0�0
1121@1Y1o1�1�1(2.2=2F2O2X2b2v23N3^3c3h3m3�3�3�3�3V4b4�4�4�4�4�4�4�4�45)555a5}5�5�5�5 664696>6q6v6{6�6�6�7�7�7�7�7�788=8B8I8�8�8�89909<9W9g9s9�9�9�9�9�9�9::u:{:�:�:�:�:�:�:�:;�;�;�;�;�;�;&<3<@<M<e<�<�<�<�<�<�<�<�<$=;=}=�=�=>B>I>[>b>�>�>�>�>�>!?)?f?o?�?�?�?   �  �   %0-0X0�0�0�0�0�0�012x2�2�2�2�23)373D3�3�3�3�4�4�4%515<6|6�6�6�6�67;7o7�7�7�7�7�78?8e8�8�8�87:�:;+;�;(<-<?<b<�<�<�<=2=d=v=�=�=�=�=>>>s>�>�>	??D?O?[?�?�?�?�?�? �  �   000"0,0T0�0�0�0�0�0"1,1Q1�12g2�2)3k3�3�4$5+5T5X5\5`5d56G6l6�6�9�9':3:�:�:�:�:�:G;|;�;�;�;�;�;�;<<F<�<�<%=,=X=i=�=�=�=c>l>�>�> �  �   �0�0�0�0�0�0�0 1)1O1m1t1x1|1�1�1�1�1�1�1�1�1�1�1R2]2x22�2�2�2�2�2	33333 3$3(3,3v3|3�3�3�3�4�4�4�4�5�5�5666�6�6�6�6�6I7R7[7c7x7}7�7�7�7�7�7848�8�8�8�8�8
9�9�9�9L:P:T:X:\:`:�:�:�:�:	;8;G;]<f<�<�<�<g=x?�?     �   �0
22=2B2G2l2u2�2�2�2�2�233!3J3S3}3�3�3�4�4�45�6�677#7(7,707Y77�7�7�7�7�7�7�7�7�7
88888�8�8�8�8�8�8�8�8999@9D9H9L9P9T9X9\9�9�9�9�9�9O<X<�=�=V>b>?�?     �0�0�0�0�0 1111;1G1N1x1�1�1�1�1�1222/292S2X2]2g2n2s2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�23_3j3q3�3�3�3�3�3!4*4T4Y4^4�4�4�4�45"5'5�5�5�5�56-62676�6�6�677A7F7K7�7�7*838]8b8g8�8�899X9a9�9�9�9::�:�:�:;$;N;S;X;�;�;Q<Z<�<�<�<�<�<=#=M=R=W=�=�=>:>C>m>r>w>�>�>r?~?�?�?�?     8  �0�0�0�0�0�0�0111$11161<1�1�1�1�1�122:2F2R2W2\2�2�2�2�2�2�2�2�2333"33�3�3�3�3�3�34-42474�4�4�4�4�4�4�4	55D5�5O6t6�6�6�6�6�677/74797�7�7�7�78�8�8�8�8�89%9@9M9R9X9e9j9p9�9�9�9":':,:1:d:p:|:�:�:�:�:�:�:;
;;;=;B;G;L;�;�;�;�;<"<'<,<W<\<a<�<�<�<�<�<�<�<='=Y=�=d>�>�>�>�>�>#?*?9?Y?^?c?�?�?   0 �   0!0+0=0G0g0l0q0�0�01H1T1Z1o1y1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2.252>2E2�2�2�2�2�2�2�2�2X3a3�3�3�3�3�3444C4L4v4{4�4x677�7�7�7�:;;�;�;�; @ �   g2�2�2�2�2373V3u3�3�3�3�34/4N4m4�4�56=6�67E7t7�8 9?9�9�9�9�9�9:":L:Q:V:r;~;�;�;�;�;�;+<0<5<^<�<�<�<�<(=-=2=p=w=�=�=">'>,>�>�>�>�>�>?C?K?�? P 4   )010�0�0�0�0�01
12224282P2U2b24/4846:Y: ` X   �0�0q1}1�1�1�1F2q3x3�4�4�5�5�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;X;\;`;�;�;�;�< p �   i1�2�2�2�2 33
33W3\3a3f3�3�3�3�3�7�7�728U8^8�8�8�8�8�8�89!9&9b9�9�9I:U:�:�:�:�:;;;a;�;�;�;�;�;�;
<<H<M<R<�<�<�<@=�=�=�=�=�=�=&>/>d>i>n>�>�>?!?F?�?�?�?�? � �   	0.0�0�0u1�1�1�122J2�2�23$4.4X4t5~5�5�6�6%7/7J7�7�7�7 88�8�8�8�8k9�9�9�9�9�9�9::!:-:6:D:M:[:a:j:x:�:�:�:�:�:;;:;L;m;~;�;�;�;�;'<8<A<]<{<�<�<�<=!=&=V=a=�=�=�=>	>�>�>�>�>�>c?�?�?�? � �   0
00�01,11161�1"23�3D4P4}4�4�4�4�4F5R55�5�5�56�6�6�6�677 7�7�7888a8i8�8�8�8�8�8V9]9�9�9�9�9�9�9d:k:�:�:�:�:�:�:<;D;<<><C<H<m<v<�<�<�<�<�<.=7=a=f=k=�=�=�=�=�=�>�>�>�>�>i?�?�?�?�?�? � �   1�1�172�3�4�45"5'5f5n5�5�5666y6�67
7D7P7}7�7�7?8K8x8}8�8�8�8�8�89�:�:�:�:�:";.;[;`;e;�;�;�;a<�<�<.=:=g=l=q=�=�=�>�>�>�>�>?&?P?U?Z?�?�?�?�?   � 8   000^0g0�0�0�0n1z1�1�1�1 5-5:8^8�8�;�;�;�=�=�= � p   �0�0�0H3M3_3X4]4o46(6}6�6L7�7�7�7�7�7~8�8�8�8*969f9k9p9�9�9�9�9�9�:�:;*;Z;_;d;�; <,<\<a<f<==%>,>`?g? � �   >0	1o12"2R2W2\273�3�3�3�34&4�9�9�9�9�9L:P:T:X:\:`:d:h:l:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�: ;;;;;;i=�>�>?!?H?T?`?v?�? � �   
00N0S0X0~0�0�0�0�0�01(1-1?1d1�1�1�172B2X2f2�2�233�3s4�4�4�4A5O5^5t5�5�5�5�5X7]7o7�7�7�7�78/8Y8m8�89u9�9�9�9�9�9	:9:>:C:�:!;k;w;�;�;�;�;�<�<�=�=�>�>�? � �   �0	1�1�1�1�1�1�2^3e3�3�3�3�3X9d9�9�9�9�9�9�9�9�9 :::::::: :8:<:@:D:H:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:)<�<�<�< =�=�=�?�?   �   0^0�0"1�1�1 22 2(2/2H2M2_2�2�2�2�2�2r3{3�3�3�3X4]4o4�4�4�4�455,5D5M5w5|5�5�5�5�56#66�688�8�8�9�9�9!:D:M:�:�:�:�:�:�:;;;K;�;�;�;<=<P<u<�<�<&=J=z=�=�=�=!>o>    �   $1(1,181<1@1D1H1T1X1\1�1�1�1 22222222 2$2(2,2024282<2@2d2h2�2�2�2`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3x6|6�6�6�6�6�8�8�8�8�8L:P:T:X:\:      �?�? 0 <   ::::$:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�?�?�?   @ �   �3�3�3�>�>�>�>�>�>�>�>�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   P 8    00000000 0$0(0,0004080<0@0D0H0L0P0T0X0   � �   �5�5�5�5�8�8�8�; <<<(<,<0<4<<<T<X<p<�<�<�<�<�<�<�<�<�<�<�<�<�<===0=@=D=T=X=\=d=|=�=�=�=�=�=�=�= > ><>@>`>|>�>�>�>�>�>�>??0?P?p?�?�?�?�?   � |   000L0P0p0�0�0�0�0�0114181T1X1x1�1�1�1�1�1�1202P2X2`2h2l2t2�2�2�2�2�2�2�2�2�233,303L3P3`3�3�3�3�3�34404P4p4   � `  0080T01111 1$1(1,10141D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�12222$2t2x2�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4D4H4L4P4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 555h5x5�5�5�5�5�5�5�5�5�5:�<�<�<�<�<�<�<�<�<�<�<�<�<====== =$=(=,=0=4=h=p=�?   �    0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          