MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       ���om��om��om�}!���om����om��ǔ�om�����om��ol��om��Ɣ�om�����om����om�Rich�om�                        PE  L нQ        � !
    �      P5                              @    ��  @                   � L   �� (    � �                     �                                  �� @                                         .text   �                        `.rdata  \�      �                @  @.data   �5   �     �             @  �.rsrc   �   �     �             @  @.reloc  `>      @   �             @  B                                                                                                                                                                                                                                                                                                                                                U���,  SVWQ�������K   ������Y�M�j hp!�������   ������P�  ���������1  �E�E�E�P�M��  ������P�M��   P�*  ����������   �M��  �M��L  �E�}� u��   R��P�� �/!  XZ_^[��,  ;���   ��]� �I    � ����   � fn �������������U����   SVWQ��4����3   ������Y�M���E�P� ��Q�B�Ѓ�;��   ��EPj��MQ�U�R� ��H�Q�҃�;��X   �E�_^[���   ;��E   ��]� ���������������U����   SVWQ��4����3   ������Y�M���E�P� ��Q�B�Ѓ�;���  _^[���   ;���  ��]������������U����   SVWQ��4����3   ������Y�M�� ����   ��M��B(��;��  _^[���   ;��  ��]��������������U���0  SVW�������L   ������h�!� ���Ph$�j��  �������������� t�������  �������
ǅ����    j h�!������7���j h�!��,����%���������Qj h�!����������P�����R������i  ���r   Pj ��,���PhJ �  ��������������z  �������O�����,����D���������9���������_^[��0  ;��S  ��]����������������U����   SVWQ��4����3   ������Y�M��E�� _^[��]��U����   SVWQ��4����3   ������Y�M��M��   �E�� "�E�_^[���   ;���  ��]������U����   SVWQ��4����3   ������Y�M��M��   �E��t�E�P�  ���E�_^[���   ;��n  ��]� ��������U����   SVWQ��4����3   ������Y�M��M��e  �E�� D"�E�_^[���   ;��  ��]������U����   SVWQ��4����3   ������Y�M��M��   _^[���   ;���  ��]��U����   SVWQ��4����3   ������Y�M��M��u  _^[���   ;��  ��]��U����   SVWQ��4����3   ������Y�M��M������E��t�E�P�d  ���E�_^[���   ;��>  ��]� ��������U����   SVW��@����0   ������������u3���   _^[���   ;���  ��]�������������U����   SVW��@����0   ������_^[��]������������U����   SVW��@����0   ������3�_^[��]����������U����   SVWQ��4����3   ������Y�M��M��5   ��E�P� ��Q$�BD�Ѓ�;��7  �E�_^[���   ;��$  ��]�U����   SVWQ��4����3   ������Y�M���E�P� ��Q�B�Ѓ�;���  �E�_^[���   ;���  ��]���������U����   SVWQ��4����3   ������Y�M��M��u�����E�P� ��Q$�BD�Ѓ�;��w  ��EP�M�Q� ��B$�H�у�;��U  �E�_^[���   ;��B  ��]� ������������U����   SVWQ��4����3   ������Y�M��M��������E�P� ��Q$�BD�Ѓ�;���  ��E�P�MQ� ��B$�HL�у�;���  �E�_^[���   ;��  ��]� ������������U����   SVWQ��4����3   ������Y�M���E�P� ��Q$�BH�Ѓ�;��_  �M��'���_^[���   ;��G  ��]����U����   SVWQ������9   ������Y�M���E�P�� ���Q� ��B$�H�у�;���  P�M�/   �� ��������E_^[���   ;���  ��]� �����������U����   SVWQ��4����3   ������Y�M���E�P� ��Q�B�Ѓ�;��  ��E�P�MQ� ��B�H�у�;��]  �E�_^[���   ;��J  ��]� ����U����   SVWQ������<   ������Y�M���E�P�����Q� ��B$�H �у�;���  P�M����������D����E_^[���   ;���  ��]� �����������U����   SVWQ��4����3   ������Y�M���E�P�MQ� ��B$�HL�у�;��{  �E�_^[���   ;��h  ��]� ��U����   SVW������9   ������EP�M�������EP�M�Q� ��B$�H@�у�;��  �E�P�M������M��`����ER��P�� �  XZ_^[���   ;���  ��]�   � ����   � fn �U���$  SVW�������I   ������ǅ8���    �=� t!������P���=�����8����������������������8���������������������������R�M������8�����t��8����������~�����8�����t��8�����������a����E_^[��$  ;���  ��]�����������U����   SVW��@����0   �������EP�MQ� ��B�H@�у�;��  _^[���   ;��  ��]�������������U����   SVW��@����0   �������EP�MQ�UR�EP�MQh�.  � ��B���   �у�;��,  _^[���   ;��  ��]���������U����   SVW��@����0   �������EP� ��Q�B�Ѓ�;���  _^[���   ;���  ��]�U����   SVW��@����0   �������EP�MQ� ��B���   �у�;��}  _^[���   ;��m  ��]����������U����   SVWQ������<   ������Y�M���E�P�M�Q�U�R�E�P� ��Q���   �Ѓ�;��  ��u3���E�R��P�� �&  XZ_^[���   ;���  ��]�   � ����    ����    ����   � data sub_id main_id U����   SVWQ��4����3   ������Y�M���E�P� ����   ��Ѓ�;��]  _^[���   ;��M  ��]����������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E�_^[��]�U����   SVWQ��4����3   ������Y�M��E��M��E��@    �E��@    �E�_^[��]� �����U���  SVWQ�������E   ������Y�M��M��E���h�  ������u���P�������	  j �E�P������Q�M��d  ������������������\  ��������t�M�����M������E��M��T   P�M������M��c����ER��P�� �!  XZ_^[��  ;���  ��]� �   � ����   � dat U����   SVWQ��4����3   ������Y�M���E�P� ����   �BL�Ѓ�;��|  _^[���   ;��l  ��]���������U����   SVW��@����0   ������j0j �)   ��P�EP�L�����_^[���   ;��  ��]������U����   SVW��@����0   ������EE_^[��]������U����   SVW��@����0   ������E� �� �� _^[��]�������������U����   SVW��@����0   ������EP�M���   Q�UR�{  ��_^[���   ;��X  ��]�����U���  SVWQ��\����i   ������Y�M��h  �M���E��8 u��   �EP��l����G���j h�"�������5���P�������)���j j���l���Q������R������P������P������Q�[�����P�����R�K�����P�E���  ������؈�c�����������������������������������������������������'�����l���������c�����t�E�P��  ���E�_^[�Ĥ  ;��"  ��]� ������������U����   SVWQ��4����3   ������Y�M��E�P�t  ��_^[���   ;���  ��]��������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   @_^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��   _^[��]� ���������������U����   SVWQ��4����3   ������Y�M��M�u����E_^[���   ;��  ��]� ������������U����   SVWQ��4����3   ������Y�M�3�_^[��]� ��U����   SVWQ��4����3   ������Y�M�3�_^[��]� ��U���  SVW��x����b   ������} u3��   j h�   ��<���P�2������E��\����E��|����E�E��E��<���ǅ@����( �E��% �E��% �E��% �E��% �E�& �E��% �E��% �E� & h�   ��<���P�MQ�URj�������R��P��% �o  XZ_^[�Ĉ  ;��-  ��]Ð   �% <����   �% np ̋�`����������̋�` ����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`����������̋�`�����������U����   SVW��4����3   ������}s�E   �E��P��  ���E��}� u3��:�} t�E��Pj �M�Q�A  ���E�� �����E����E���   �E�_^[���   ;���
  ��]������������U����   SVW��4����3   ������} tF�E�E��=� t�E�x��u�E��P�h  �����E�P� ��Q��Ѓ�;��
  _^[���   ;��v
  ��]���U����   SVW��<����1   ������= � tI�}sǅ<���   �	�E��<�����MQ�UR��<���P� ��Q���   �Ѓ�;��
  �j�EP�e�����_^[���   ;���	  ��]���������������U����   SVWQ��4����3   ������Y�M��E�� �"�E�_^[��]�����������U����   SVWQ��4����3   ������Y�M��M��5   �E��t�E�P�d������E�_^[���   ;��>	  ��]� ��������U����   SVWQ��4����3   ������Y�M��E�� �"_^[��]��������������U����   SVWQ������=   ������Y�M��E��E�}� tM�E쉅 ����� ������������� t%��j��������������;��  ������
ǅ���    �E�    _^[���   ;��]  ��]����������U����   SVW��<����1   ������E��<�����<���t��E���E���   _^[��]� U����   SVW������:   ������E�����������������������q  ������$�|+ �   �]  �������=���   �EP������=�.  }
������&  �} u
������  h�"�P���Ph$�j��������� ����� ��� t�� �������������
ǅ���    ��������=� t�EP���2����   �   �EP�MQ�+�������u����   �   �|�����u������u\������  �=� t?����8�����8�����,�����,��� tj��,����_   ������
ǅ���    ��    �   ����_^[���   ;��9  ��]Ð
* �* �*  * d+ �* ������������U����   SVWQ��4����3   ������Y�M��M��E����E��t�E�P��������E�_^[���   ;��  ��]� ��������U����   SVW��@����0   ������h ��EPhD ��  ��_^[���   ;��l  ��]���������U����   SVWQ��(����6   ������Y�M�j\�������E�}� t	�E�x\ u�$��E�P�M�Q\�҃�;��  �EP�M��   �E�_^[���   ;���  ��]� ��U����   SVWQ��(����6   ������Y�M�j`�������E�}� t	�E�x` u���E�P�M�Q`�҃�;��  _^[���   ;��w  ��]����U����   SVWQ��(����6   ������Y�M�jd�������E�}� t	�E�xd u���EP�M�Q�U�Bd�Ѓ�;��  _^[���   ;��  ��]� �������������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR� ����   �M��B��;��  _^[���   ;��  ��]� ���������������U����   SVWQ��4����3   ������Y�M��E��     �E��@    �E��@    �E��@    �E�_^[��]�������������U����   SVWQ��4����3   ������Y�M��M��   _^[���   ;���  ��]��U����   SVWQ������:   ������Y�M��E��x t�   �E��8 t)��E��Q� ��B<�H�у�;��  �E��     �E��x tS�E��x t@�E��H��,�����,����� ����� ��� tj�� ����.���������
ǅ���    �E��@    _^[���   ;��  ��]���������������U����   SVW��@����0   ������������_^[���   ;���  ��]�����U����   SVW��@����0   ������ ��H����;��  _^[���   ;��}  ��]����������U����   SVW��@����0   �������E�Q� ��B�H�у�;��2  �E�     _^[���   ;��  ��]������U����   SVWQ��4����3   ������Y�M���EP�MQ�UR�E�P� ��Q�B�Ѓ�;���   _^[���   ;��   ��]� �������������U����   SVW��(����6   ������} t�E�8 t�E� �Pj�EP�������E��}� u3��5�M�������E�}� u3�� �} t�E�M��E�M;H~3���E�_^[���   ;��   ��]����������u�U��� PRSVW�Ej P�w  ��_^[ZX��]�����������̋�U��QSVW3���ى}�9>~H���$    ��F�8�|�����u�T8с<����t�L8�UQR��  ���E�@���E�;|�_^[��]�����������̀=%� uj jj j j �%���  P�{  ����������jjj j j �  ���������������̋�U��Q�M��E�� �"�M�Q�  ����]��������������̋�U��Q�M��M������E��t�M�Q��������E���]� �̋�U��Q�M��E���	P�M��	Q�d  ���������]� ���̋�U��j�h(�h � d�    P���SVW�t�1E�3�P�E�d�    �}��   �/N  ��u3��  ��  ��u�VN  3��  �M  � ����L  �,��A  ��}��  �"N  3��i  ��G  ��|�=F  ��|j ��;  ����t�E  �  ��M  3��3  j�n;  ���(����(��  �} um�=(� ~X�(����(��E�    �=�� u�<  �!E  �,  �M  �E������   ��} u�=���t�  ��3��   �   �}��   �  h�   h�"jh  j�/  ���E�}� tV�U�R���P�\�Q� �Ѕ�t%j �U�R��  ���  �M��U��B�����j�E�P��#  ��3���3����}u
j ��  ���   �M�d�    Y_^[��]� �������������̋�U��}u��N  �EP�MQ�UR�   ��]� �������̋�U��j�hH�h � d�    P���SVW�t�1E�3�P�E�d�    �e��E�   �} u�=(� u3��N  �E�    �}t�}uT�=�" t�EP�MQ�UR��"�E�}� t�EP�MQ�UR�����E�}� u�E�    �E������E���   �EP�MQ�UR�����E�}u=�}� u7�EPj �MQ������URj �EP�����=�" t�MQj �UR��"�} t�}u@�EP�MQ�UR������u�E�    �}� t�=�" t�EP�MQ�UR��"�E��E������8�E���U��E�P�M�Q�N  ��Ëe��E�    �E������E��
�E������E�M�d�    Y_^[��]��������������̋�U���   �} t�;P  ��]�������̋�U��� �� ���� ��p� ��Ї ���� ��� ��P� ��� � �Ј �$��� ]������;t�u����g  ̃=�� �Ct  ���\$�D$%�  =�  u�<$f�$f��f���d$�t  � �~D$f(0#f(�f(�fs�4f~�fT`#f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�Fh  ���D$��~D$f��f(�f��=�  |!=2  �fT #�\�f�L$�D$����f�P#fVP#fT@#f�\$�D$���������������̃=�� t-U�������$�,$�Ã=�� t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������̋T$�L$��ti3��D$��u���   r�=�� t�s  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$������̋�U��Qj j j���P�MQ�e  ���E��E���]��������̋�U��j�EP�`  ��]������������W�|$�n��$    ���L$W��   t�����t=��   u�������~Ѓ��3�� �t�A���t#��t�  � t�   �t�͍y���y���y���y��L$��   t�����tf�����   u���������~�Ѓ��3��� �t��t4��t'��  � t��   �t�ǉ�D$_�f��D$�G _�f��D$_È�D$_��������̀�@s�� s����Ë���������������������������̺p#�!�  �p#霁  ���������z�����������������̋�U��j�hh�h � d�    P���SVW�t�1E�3�P�E�d�    �)8  �E�    �EP�9   ���E��E������   �� 8  ËE�M�d�    Y_^[��]����������̋�U������P� �E����Q� �E��U�;U�r�E�+E�����s3���   j�M�Q�!  ���E�U�+U���9U���   �}�   s�E�E���E�   �M�M�M�U�;U�r"j}h�#j�E�P�M�Q�*  ���E��}� u:�U���U�E�;E�r%h�   h�#j�M�Q�U�R��  ���E��}� u3��Q�E�+E����M����U��E��E��M�Q� ����UR� �M���U����U��E�P� ����E��]���������������̋�U��EP�"���������؃�]����̋�U��Qh�   h�#jjj ��  ���E��E�P� ����������}� u�   ��U��    3���]��������̋�U��E��w$�������&���tRP�EQP�4   ��]ú�#R�   P�E�   QP�   ��]���������������̋�U���@  �t�3ŉE��ES�]VW�}S������������ǅ����    �C  ����������uS�   ���������5 j j j�Wj h��  ��=   s&P������Qj�Wj h��  �օ�t�������������
ǅ�����'h  �p  ����������t%���������&PSQW��  �����"  2��������� ������u���  ��t� ����   h  ������R������Ph  ������Q���S�;�  ����t-������������RWh�'������P�EQ������RP���   �= j j h
  ������Qj�������Rj h��  �h'�ׅ�t������j j h
  ������Pj�������Qj h��  �T'�ׅ�t������������������������R�UPh4'VQSR����������u̋M�_^3�[�#�����]���������������̋�U��j�h��h � d�    P��$SVW�t�1E�3�P�E�d�    �e�3��E��E�  �M�MЍU�UԉE��M�QjPh�m@� �	�   Ëe��E������E�M�d�    Y_^[��]������̋�U��j�h��h � d�    P��$SVW�t�1E�3�P�E�d�    �e�3��E��E�  �M�MЋU�UԋM�M؍U�U܋M�M��E��U�RjPh�m@� �	�   Ëe��E������E�M�d�    Y_^[��]����̋�U���  �t�3ŉE��=����E�������E��   �8 SV��   �ȍq���A��u�+΃�-��   w{������3ɍd$ ���&������A��u�Њ@��u�W������+�O�OG��u��������ȃ���&�Ȋ@��u�������+���O�OG��u������ȃ��_��,(���������SjPQ�������^[�M�3��������]����̋�U��M�H��H��D�    ]�̡D�����������̡H�����������̋�U��0� ]����̋�U��j�hȞh � d�    P���SVW�t�1E�3�P�E�d�    j�ǒ  ���E�    �E�x ��   �P��M��E�L���U��U�}� tV�E�M�;Qu�E��M�Q�P�E�P�������/�M�M��U�z uh�)j jXh()j�7�  ����u�랋M�QR�`������E�@    �E������   �j�N�  ��ËM�d�    Y_^[��]��������̋�U��} u��EP�MQ�UR�EP�MQ�J�  ]��������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t�����������̋�U��j � ]�̋�U���( ]� ̋�U��Q���P�, �E��}� u �X�Q� �E��U�R���P�0 �E���]��������������̋�U���h,*�8 �E��}� u��  3���  h *�E�P�  �T�h*�M�Q�  �X�h*�U�R�  �\�h *�E�P�  �`��=T� t�=X� t�=\� t	�=`� u,�T� E �, �X��0 �\��4 �`��( ����=���t�X�Q���R�0 ��u3���   �.  �T�P� �T��X�Q� �X��\�R� �\��`�P� �`��Ռ  ��u�   3��   h J �T�Q� �У���=���u	�~   3��rh  h�)jh  j��
  ���E��}� t�U�R���P�\�Q� �Ѕ�u	�4   3��(j �U�R�   ���  �M���U��B�����   ��]����̋�U��=���t���P�`�Q� ����������=���t���R�4 ��������^�  ]������������̋�U��j�h�h � d�    P���SVW�t�1E�3�P�E�d�    h,*�8 �E�E�@\�:�M�A    �U�B   �E�@p   �MƁ�   C�UƂK  C�E�@h�j�Ӎ  ���E�    �M�QhR�< �E������   �j��  ���j蜍  ���E�   �E�M�Hl�U�zl u�E�ص�Hl�U�BlP�ȕ  ���E������   �j萍  ��ËM�d�    Y_^[��]����������̋�U����D �E����P�����ЉE��}� u}j h�  h�)jh  j�  ���E��}� tW�M�Q���R�\�P� �Ѕ�t%j �M�Q�[������  �U���E��@�����j�M�Q�6  ���E�    �U�R�@ �E���]�����������̋�U��Q�5����E��}� u
j�&  ���E���]�����������̋�U��j�h�h � d�    P���SVW�t�1E�3�P�E�d�    �E�E܃}� ��  �M܃y$ tj�U܋B$P�  ���M܃y, tj�U܋B,P�m  ���M܃y4 tj�U܋B4P�S  ���M܃y< tj�U܋B<P�9  ���M܃y@ tj�U܋B@P�  ���M܃yD tj�U܋BDP�  ���M܃yH tj�U܋BHP��  ���M܁y\�:tj�U܋B\P��  ��j�$�  ���E�    �M܋Qh�U��}� t%�E�P�H ��u�}��tj�M�Q�  ���E������   �j��  ���j�Ɗ  ���E�   �U܋Bl�E�}� t4�M�Q�$�  ���U�;صt�}� �t�E�8 u�M�Q�,�  ���E������   �j褊  ���j�U�R��  ���M�d�    Y_^[��]� �������������̋�U��=���tO�} u)���P�, ��t���Q���R�, �ЉEj ���P�\�Q� �ЋUR�����=���tj ���P�0 ]����������̋�U��Q�EP�MQ�UR���P�MQ�   ���E��E���]��̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�4   ���E��}� u�}� t譥  ��t
褥  �M���E���]��������̋�U��Q�EP�MQ�UR�EP�MQ�a   ���E��}� t�E��?�} u�} t	�U�   �E��%�EP譥  ����u�} t	�M�   3��뗋�]�������������̋�U��j�h8�h � d�    P���SVW�t�1E�3�P�E�d�    �E�    �E�    j�Y�  ���E�    �=�� vU�����9l�u6�a  ��u!h�+j h  h8+j��  ����u��l�    ��l����l�����E؃=���t�M�;��u̃=p� tu�UR�EP�M�Q�UR�EPj j�p�����uP�} t%�MQ�URh +j j j j �|  ����u�� h�*hh"j j j j ��{  ����u��D  �U����  ��t�����u�E�   �}�v3�MQh�*j j j j�{  ����u̃} t	�E�    ��  �M����  ��t:�}t4�U����  ��t&�}t h�*hh"j j j j�?{  ����u̋M��$�MԋU�R��  ���E܃}� u�} t	�E�    �r  ���������}� tI�U��    �E��@    �M��A    �U��B�����E܋M�H�U��B   �E��@    �   ���+d�;Mv�d�U�d��
�d������|�E�|��|�;p�v�|��p��=t� t�t��M܉H�	�U܉h��E܋t���U��B    �E܋M�H�U܋E�B�M܋U�Q�E܋M�H�U܋E؉B�M܉t�j���R�E܃�P�������j���Q�U�E܍L Q�������UR���P�M܃� Q�������U܃� �U��E������   �j�=�  ��ËE��M�d�    Y_^[��]����̋�U��Q�} v�����3��u;Es�0�  �    3��K�E�E�E�MQ�UR�EP�MQ���R�EP�l������E��}� t�MQj �U�R��������E���]�������̋�U����E�    �E�P�MQ�UR�EP�MQ�UR�T������E��}� u�}� t荠  ��t
脠  �M���E���]��������̋�U��j�hX�h � d�    P���SVW�t�1E�3�P�E�d�    j�ǃ  ���E�    j�EP�MQ�UR�EP�MQ�B   ���E��E������   �j�ǃ  ��ËE�M�d�    Y_^[��]��������������̋�U����E�    �E��M��} u�UR�EP�MQ�U�R�~������  �} t�}� u�EP�MQ�  ��3��  �=�� vV�����9l�u6�  ��u!h�+j h�  h8+j�{  ����u��l�    ��l����l�����U�=���t�E�;��u̃=p� ty�MQ�UR�E�P�MQ�U�R�EPj�p�����uR�} t%�MQ�URh�.j j j j �v  ����u�� h|.hh"j j j j �v  ����u�3��  �}��v`�} t)�UR�EP�M�Qh8.j j j j�Zv  �� ��u���E�Ph�*j j j j�9v  ����u���  �    3��3  �}th�U����  ��tZ�E%��  ��tM�} t%�MQ�URh�-j j j j��u  ����u�� h�*hh"j j j j�u  ����u��Qj���R�E�����P�  ����t1�MQh�-j j j j�zu  ����u��\�  �    3��t  �EP��  ����u!hP-j h  h8+j�y  ����u̋U�� �U�E�xu�E�   �}� t8�M�y����u	�U�z t!h�,j h#  h8+j�Ry  ����u��d�M�Q����  ��u�E%��  ��u�E   �M�d�;Qs1�EPh�,j j j j�t  ����u��p�  �    3��  �} t%�U���$R�E�P荞  ���E��}� u3��_  �#�M���$Q�U�R��  ���E��}� u3��:  3�u����������}� u|�=d��s9�U�d�+B�d����+d�;M�v�d�U��d��
�d������E��|�+H�|��|�U��|��|�;p�v�|��p��U��� �U�E��M�;Hv$�U��E�+BP���Q�U��E�BP�[�����j���Q�U�U�R�B������}� u�E��M�H�U��E�B�M��U�Q�E��M��H�} u/�} u�U�;U�t!h(,j h�  h8+j�Yw  ����u̋M�;M�t�}� t�E���   �U��: t�E���U��B�A�8�h�;M�t!h�+j h�  h8+j��v  ����u̋E��H�h��U��z t�E��H�U����7�t�;M�t!h�+j h�  h8+j�v  ����u̋E���t��=t� t�t��E��B�	�M��h��U�t���M��A    �U��t��E��]�������̋�U��j�hx�h � d�    P��SVW�t�1E�3�P�E�d�    j�'}  ���E�    �EP�MQ�0   ���E������   �j�8}  ��ËM�d�    Y_^[��]��̋�U��Q�=�� vU�����9l�u6��  ��u!h�+j h  h8+j�u  ����u��l�    ��l����l��} u�l  �}uOj���P�M�����Q�B  ����t/�URh�2j j j j�p  ����u�藘  �    �  �=p� tDj j j �MQj �URj�p�����u%h�2hh"j j j j �]p  ����u���  �MQ�  ����u!hP-j h*  h8+j�t  ����u̋E�� �E��M��Q����  ��tD�E��xt;�M��Q����  ��t*�E��xt!hx2j h0  h8+j�9t  ����u̋�����m  j���P�M���Q�  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��l*Ph�1j j j j�Eo  ��(��u��<�U��� R�E��HQ�U��B%��  ��l*Qh@1j j j j�o  �� ��u�j���P�M��Q�E��L Q�Q  ������   �U��z tM�E��HQ�U��BP�M��� Q�U��BP�M��Q����  ��l*Ph�0j j j j�n  ��(��u��<�U��� R�E��HQ�U��B%��  ��l*Qh0j j j j�Mn  �� ��u̋E��xue�M��y����u	�U��z t!h�/j hi  h8+j�~r  ����u̋M��Q��$R���P�M�Q��������U�R�~  ���Q  �E��xu�}u�E   �M��Q;Ut!hT/j hw  h8+j�r  ����u̋M��|�+Q�|��������   �M��9 t�U���M��Q�P�6�h�;E�t!h(/j h�  h8+j�q  ����u̋U��B�h��M��y t�U��B�M����5�t�;E�t!h�.j h�  h8+j�\q  ����u̋U���t��M��Q��$R���P�M�Q�������U�R��|  ���(�E��@    �M��QR���P�M��� Q��������]�̋�U��j�h��h � d�    P���SVW�t�1E�3�P�E�d�    3��} ���E܃}� u!h�.j h�  h8+j�p  ����u̃}� u1� �  �    j h�  h8+h43h�.�|  ������8  �=�� vV�����9l�u6�u  ��u!h�+j h�  h8+j�p  ����u��l�    ��l����l�j��v  ���E�    �UR��  ����u!hP-j h�  h8+j�o  ����u̋M�� �M��U��B%��  ��tC�M��yt:�U��B%��  ��t*�M��yt!hx2j h�  h8+j�`o  ����u̋E��xu�}u�E   �M��Q�U��E������   �j�sv  ��ËE�M�d�    Y_^[��]����������̋�U��E�M���M��t�U�E��E���E;�t3���Ӹ   ]�������̋�U��j�h��h � d�    P���SVW�t�1E�3�P�E�d�    �����u
�   ��  j�u  ���E�    �$�  �E��}����   �}����   �M��MЋUЃ��UЃ}���   �E��$��d h�5hh"j j j j �i  ����u��   hd5hh"j j j j �~i  ����u��dh@5hh"j j j j �\i  ����u��Bh5hh"j j j j �:i  ����u�� h�4hh"j j j j �i  ����u��E�    ��  �E�   �t��E���M��U�}� ��  �E�   �E�H����  ��t#�U�zt�E�H����  ��t	�U�zu�E�H����  ��l*�U���E��4j���P�M��Q���������uz�U�z t=�E�HQ�U�BP�M�� Q�U�BP�M�Qh�1j j j j �.h  ��(��u��-�E�� P�M�QR�E�Ph@1j j j j ��g  �� ��u��E�    j���R�E�H�U�D
 P�B�������uz�M�y t=�U�BP�M�QR�E�� P�M�QR�E�Ph�0j j j j �g  ��(��u��-�U�� R�E�HQ�U�Rh0j j j j �ag  �� ��u��E�    �M�y ��   �U�BP���Q�U�� R��������ud�E�x t2�M�QR�E�HQ�U�� RhH4j j j j ��f  �� ��u��"�M�� Qh�3j j j j ��f  ����u��E�    �}� uz�E�x t=�M�QR�E�HQ�U�BP�M�� Q�U�Rhx3j j j j �}f  ��(��u��-�M�QR�E�� P�M�QhL3j j j j �Nf  �� ��u��E�    �G����E������   �j��q  ��ËE܋M�d�    Y_^[��]ÍI oa Ma +a a �������̋�U��j�h؟h � d�    P���SVW�t�1E�3�P�E�d�    ����E�}�t�M����  ���t	�E�    ��E�   �U܉U��}� u!h�5j hy  h8+j��i  ����u̃}� u0�J�  �    j hy  h8+h�5h�5��u  ������sj�p  ���E�    ����M�}�t7�U��t���   ��E��%��  ����l�    �M����E������   �j�p  ��ËE�M�d�    Y_^[��]����������̋�U��3��} ��]Ë�U��} u3��1j j �E�� P���������u3���M�� Qj ���R�L ]��������������̋�U��j�h��h � d�    P���SVW�t�1E�3�P�E�d�    3��} ���E܃}� u!h�7j h�  h8+j�Th  ����u̃}� u.���  �    j h�  h8+h�7h�7�Ot  ���m  j� o  ���E�    �U�t���E�    �	�M���M�}�}�U�E�D�    �M�U�D�    �ӡt��E���M���U��}� ��   �E��H����  |f�U��B%��  ��}V�M��Q����  �E�L����U��B%��  �U�L��E��H����  �U�D��M�A�U��J����  �U�D��W�E��x t/�M��QR�E��HQ�U�Rht7j j j j �b  �� ��u���M�QhP7j j j j �xb  ����u������E�p��H,�U�d��B0�E������   �j��m  ��ËM�d�    Y_^[��]��������̋�U����E�    �E�P�M��%   �M��-  P�MQ�3  ���M���   ��]����̋�U��Q�M��E��@ �} ��   ������M��A�U��B�M��Pl��E��H�U��Ah�B�M��;صt�E��H�Qp#t�u
�{  �M���U��B;�t�M��Q�Bp#t�u�{  �M��A�U��B�Hp��u�U��B�Hp���U��B�Hp�M��A��U��J�U���J�E���]� ������̋�U��Q�M��E��H��t�U��B�Hp����U��B�Hp��]���̋�U��Q�M��E���]Ë�U��j�h�h � d�    P���SVW�t�1E�3�P�E�d�    �E�    j� l  ���E�    h�8hh"j j j j �_`  ����u̃} t�M��U�t��E���M��U�}� �(  �E�;E��  �M�Q����  ��t)�E�H����  t�U�B%��  ��u�����u��  �U�z twj j�E�HQ�(�������tj�U�BP�P ��t$�M�QRh�8j j j j �_  ����u��)�M�QR�E�HQh�8j j j j �j_  ����u̋E�HQh�8j j j j �H_  ����u̋E�H����  ����   �U�BP�M�Q������  R�E�� Phd8j j j j ��^  �� ��u̃=x� t,j�U�� R�P ��u�E�HQ�U�� R�x�����E�P�MQ��   ���   �U�zu;�E�HQ�U�� Rh<8j j j j �~^  ����u̋M�Q�UR�   ���Z�E�H����  ��uI�U�BP�M�Q������  R�E�� Ph8j j j j �"^  �� ��u̋U�R�EP�\   ��������E������   �j�i  ���h�7hh"j j j j ��]  ����u̋M�d�    Y_^[��]���������̋�U���t�t�3ŉE��EP�M������E�    �	�M����M��U�z}�E�H�M���E�   �U�;U��  �EE��H �M��M��u�����t3�M��i�������   ~ �M��V���PhW  �E�P�։  ���E��hW  �M�Q�M��,���P��  ���E��}� t	�U��U���E�    �E��M��L�軄  ��U�豄  �     �E�PhX(�M�k��1   +�R�E�k��L�Q��  ����}*j h	  h8+h�8h�8j"j�]�  �R�U   �� �M�  �M��������U��D� �E�P�M�Qh�8j j j j �1\  ����u̍M�� ����M�3��&�����]��̋�U��} t�E;Et�M;Mt�E��U$R�E P�MQ�UR�EP��l  �E]��̋�U���8�t�3ŉE��E�P�u������}� u�}� u�����t7�}� t1h$9hh"j j j j �~[  ����u�j �N������   �3��M�3��h�����]����̋�U��Q����E��E���]�����������̋�U�졀�]����̋�U��Q�=# th#�7�  ����t�EP�#���/  hL!h4!�?  ���E��}� t�E��Ghp� �������h0!h !��  ���=�� th���̌  ����tj jj ���3���]���̋�U��j j�EP�  ��]���������̋�U��jj j �  ��]�����������̋�U���Q  �EP�-R  ��h�   ����]��������������̋�U��Q����E��	�M����M��}� t�U��: tj�E��Q���������j���R����������    ����E��	�M����M��}� t�U��: tj�E��Q��������j���R���������    j���P������j���Q�p�����j���R� P�X��������    ���    �l��������P�H ��u'�=��tj��Q�����������R�< ��]���������������̋�U��j�h8�h � d�    P���SVW�t�1E�3�P�E�d�    �  �E�    �=���U  ���   �E����} ��   ���Q� �E�}� ��   ���R� �E��E�    �E�EԋM؉M�   ����   �E�    �E�    �E؃��E؋M�;M�r�;����U�9u��E�;E�s�h�M؋R� �E������M؉�U܋��R� �EС��P� �E̋M�;M�u�U�;U�t�EЉEԋMԉM�ỦU��E��E��T���h`!hP!�  ��hh!hd!�  ���=�� u#j��L������� t���   �����P����E������   ��} t�   Ã} t����   �   �MQ�V   ���M�d�    Y_^[��]�̋�U���hL9�8 �E��}� th<9�E�P�  �E��}� t�MQ�U���]�̋�U��EP�������MQ�T ]���̋�U��j��a  ��]���������������̋�U��j�b  ��]���������������̋�U��Q�u����E��E�P�i~  ���M�Q�f  ���U�R�AQ  ���E�P�u�  ���M�Q虊  ���U�R�-�  ����]������̋�U��E;Es�M�9 t�U��ЋM���M��]�������̋�U��Q�E�    �E;Es#�}� u�M�9 t
�U��ЉE��M���M�ՋE���]�̋�U���p�E�P�h h�   hd9jj@j �Y������E��}� u�����  �M�������    �	�U���@�U����   9E�s^�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B$$�M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��E����  �}� ��  �M��U��E���E��M�M��M��}�   }�U��U���E�   �E��E��E�   �	�M����M����;U���   h�   hd9jj@j �6������E��}� u����E��   �M��U���������� ����	�M���@�M��U�����   9E�sP�M��A �U�������E��@
�M��A    �U��B$$��M��A$�U��B%
�E��@&
�M��A8    �U��B4 ��,����E�    ��E����E��M����M��U����U��E�;E���   �M��9���   �U��:���   �E����tv�U����u�M��R�d ��t[�E����M���������M��U��E���
�U��E���Jh�  �U���R�` ��u����`  �E��H���U��J�;����E�    �	�E����E��}��!  �M������M��U��:�t�E��8���   �M��A��}� u	�E�������U�����҃���U��E�P�\ �E��}����   �}� ��   �M�Q�d �E��}� tr�U��E���M����   ��u�U��B��@�M��A��U����   ��u�E��H���U��Jh�  �E���P�` ��u����R�M��Q���E��P��M��Q��@�E��P�M��������U��B�   �M��A��������R�X 3���]�̋�U����E�    �	�E����E��}�@}y�M��<��� tg�U������E��	�M���@�M��U�����   9E�s�M��y t�U���R�l ��j�E�����Q��������U�����    �x�����]���̋�U����=�� u�w  �E�    �,��E��}� u����e  �M����t,�E����=t	�U����U��E�P�_  ���M��T�U���juhD:jj�E���P�P������E�M����=�� u�����   �,��U��	�E�E��E��M������   �E�P�^  �����E��M����=��   j~hD:jj�E�P��������M��U�: uj���P���������    ����rj h�   h�9h�9h�9�M�Q�U�R�E�Q�A[  ��P��������U���U��B���j�,�P�Z������,�    �M��    ���   3���]����̋�U����E�    �=�� u�v  ��� h  h��j �p h����   ���=�� t������t����U���E����E�E�M�Q�U�Rj j �E�P�   ���}����?s�}��r����w�M��U���;E�s����dh�   hx:j�M��U���P�������E��}� u����8�M�Q�U�R�E��M���R�E�P�M�Q�6   ���U�������E����3���]���������̋�U��E���]�̋�U����E�     �M�   �U�U��} t�E�M��U���U�E�    �E����"u3҃}� �U��E���M�U����U��w�E����U�
�} t�E�M����E���E�M���U�E����E��M�Q�ǅ  ����t/�U����M��} t�U�E���
�U���U�E����E��M��t �}� �M����U�� t�E��	�7����M��u�U����U���} t�E�@� �E�    �M����t!�E���� t�U����	u�M����M��ߋU����u��  �} t�M�U��E���E�M����E��E�   �E�    �M����\u�E����E��M���M���U����"uH�E�3ҹ   ���u0�}� t�U��B��"u�M����M���E�    3҃}� �U��E���E�M�U���U��t$�} t�E� \�M���M�U����M��̋U����t�}� u�M���� t�E����	u�   �}� ��   �} tQ�U��P��  ����t)�M�U����M���M�U����U��E����U�
�E�M����E���E�)�M��R蘃  ����t�E����E��M����E��M����E��M����M��|����} t�U� �E���E�M����E�������} t�M�    �U���U�E����U�
��]Ë�U����E�    �x �E��}� u3���   �E��E�M����t�E���E�M����u	�E���E��؋M�+M������M�j j j j �U�R�E�Pj j � �E��}� tjJh�:j�M�Q�������E�}� u�U�R�t 3��Dj j �E�P�M�Q�U�R�E�Pj j � ��uj�M�Q��������E�    �U�R�t �E��]��������̋�V����=�s���t�Ѓ����r�^����������̋�V� ���=$�s���t�Ѓ���$�r�^����������̋�U��Q�E�   j h   j �| ����=�� u3���   ��]���������̋�U����P�� ���    ]���̋�U���0�E� �E�   �E���E��M����M�U��B3t��EԋM�Q�U�R�  ���E�H��f�   �U�U��E�E��M��U��Q�E��H�M���U�U؃}����   �E�k��MԍT�U�E�H�MЋU��E�}� ��   �U�M��y[  �E��E��}� }�E�    �   �   �}� ��   �M�9csm�u)�=�� t h����y  ����tj�UR������M����U�?[  �E��H;M�tht��U�R�M����U��6[  �E��M�H�U�R�E�P�e   ���U�M�I��Z  �����&�U��z�tht��E�P�M����������Z  �E��M߅�t�U�R�E�P�   ���E��]��������̋�U����E�8�t%�M��E��M��U�EB3E��E��M��۳���M�Q�E��M��U�EB3E��E��M�赳����]�̋�U����E�    �E�    �=t�N�@�t�t�%  ��t�t��щx��   �U�R�� �E��E�M�3M��M��� 3E�E��  3E�E��� 3E�E�U�R�� �E�3E�E�M�3M�M�}�N�@�u	�E�O�@���U��  ��u�E�G  ��E�E�M�t��U��҉x���]Ë�U��}csm�u�EP�MQ�   ����3�]����������̋�U���������E��}� u3���  �E��H\Q�UR��  ���E��}� u	�E�    �	�E��H�M�}� u3��  �}�u�U��B    �   �  �}�u����v  �E��H`�M�U��E�B`�M��y�4  �p;�U��	�E����E��p;t;9M�}�U�k��E��H\�D    �ЋU��Bd�E�M��9�  �u�U��Bd�   �   �E��8�  �u�M��Ad�   �   �U��:�  �u�E��@d�   �   �M��9�  �u�U��Bd�   �q�E��8�  �u�M��Ad�   �Z�U��:�  �u�E��@d�   �C�M��9�  �u�U��Bd�   �,�E��8� �u�M��Ad�   ��U��:� �u
�E��@d�   �M��QdRj�U���E��M�Hd��U��B    �E��HQ�U���U��E�B`�����]������̋�U��Q�E�E��M��;Ut�E����E��|;k�M9M�s�ڋ|;k�U9U�s
�E��;Mt3���E���]��������̋�U��j jh<h�;h�;h   h   j �|  ��P莼����]���������̋�U��j �EP�   ��]�����������̋�U����EP�M�������M�R�  ����et�E���E�M�R�s}  ����u�E�Q�p  ����xu	�U���U�E��M��M���������   ��U���M���M�U��E��M�U���E��E��M��E���E��u׍M�������]Ë�U��j �EP�   ��]�����������̋�U���V�EP�M�������M���t*�E�0�M����������   ��;�t�U���U�̋E��U���U����   �E���t!�U���et�M���Et�E���E�ՋM�M��U���U�E���0u�U���U��E�0�M��b�������   ��;�u	�U���U�E���E�M�U����M��E����E���t�؍M������^��]���̋�U��Q�E�������Az	�E�   ��E�    �E���]�����̋�U����} t$�EP�MQ�U�R��}  ���E�M���U��P��EP�MQ�U�R�~  ���E�M���]��������������̋�U��j �EP�MQ�UR������]���̋�U���D�t�3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P��  ��3Ƀ} ���Mă}� u!h =j h�  h�<j�5D  ����u̃}� u3�g  �    j h�  h�<h�<h =�0P  ���   �  3�;E��ىM�u!hx<j h�  h�<j��C  ����u̃}� u3�9g  �    j h�  h�<h�<hx<��O  ���   �   �}�u�E�E���M�3҃9-�E+�3Ƀ} ��+��E��U�R�E��P�M�Q�U�3��:-��E3Ƀ} ���P�!~  ���Eȃ}� t�U� �E��(�EPj �M�Q�UR�EP�MQ�UR�   ���EȋEȋM�3�舫����]����̋�U���@�E�    �E P�M��u���3Ƀ} ���M܃}� u!h =j h3  h�<j�B  ����u̃}� u@�f  �    j h3  h�<hl>h =�N  ���E�   �M�������E���  3�;E��ىM�u!hx<j h4  h�<j�&B  ����u̃}� u@�e  �    j h4  h�<hl>hx<�!N  ���E�   �M��o����E��}  3��} ����#E��	;E��ىM�u!h�=j h<  h�<j�A  ����u̃}� u@�e  � "   j h<  h�<hl>h�=�M  ���E�"   �M�������E���  �E��t'�M3҃9-��U�U�3��} ��P�M�Q�6  ���U�U��E�8-u�M��-�U����U��} ~-�E��M��Q��E����E��M���������   ��M����E�E�M��Ƀ���E��}�u�U�U���E�+E�M+ȉM�j h_  h�<hl>h@=h8=�U�R�E�P��G  ��P萵�����M����M�} t�U��E�E����E��M�Q���0��   �M�Q���U�y�E��؉E��M��-�U����U��}�d|)�E���d   ���ЋE��ʋU��
�E���d   ���U��U����U��}�
|)�E���
   ���ЋE��ʋU��
�E���
   ���U��U����U��E��M��ЋE������t �U����0uj�M��Q�U�R�  ���E�    �M�������Eċ�]������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���   �E�E��E��  �E�    �E�    �E�    �0   f�M��E�    �E�    3�f�U��E�    �E�    �E�    �E�    �EP�M��^����} }�E    3Ƀ} ���M��}� u!h =j h�  h�<j�w>  ����u̃}� u@��a  �    j h�  h�<h�>h =�rJ  ���E�   �M�������E���  3�;E��ىM�u!hx<j h�  h�<j�>  ����u̃}� u@�na  �    j h�  h�<h�>hx<��I  ���E�   �M��K����E��g  �E�  �M��;M��ډU�u!h�>j h�  h�<j�=  ����u̃}� u@��`  � "   j h�  h�<h�>h�>�~I  ���E�"   �M�������E���  �M��Q�4�Ձ  %�  �� �E��U��}��  ��   �}� ��   �}�u�U�U��	�E���E�j �MQ�U�R�E��P�MQ�������E��}� t�U� �E��E��M��?����E��[  �M�Q��-u�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���Eje�MQ�  ���E��}� t!�U��Ҁ����p�E���M����M��U�� �E��E��M������E���  �M��Q�?赀  ���� ��|����U���|���U�t�E� -�M���M�U�0�E���E�M��ɀ����x�U�
�E���E�M��ɀ����a�у�:�U��M��Q�4�=�  %�  �� ��t�����x�����t����x���u[�E� 0�M���M�U��J���� ��l�����p�����l����p���u�E�    �E�    ��EЃ��Mԃ� �EЉM���U�1�E���E�M�M��U���U�} u�E��  ��M���������   ��M����E��P���� ��d�����h�����h��� w��d��� �p  �E�   �E�    �M܋E�U��  �E�U��E܅���   �} ~}�M��Q���� #E�#U��M���~  f�E��U���0f�U��E���9~�M�M�f�M��U�E���M���M�E�U��~  �E�U��U܃�f�U܋E���E�q����M܅���   �U��R���� #E�#U��M��p~  f�E��E�����   �M�M��U����U��E����ft�U����Fu�M��0�U����U��ًE�;E�t/�M����9u�E���U��D�M����U�����M����U����U��E�����U��
�	�E���E�} ~�M�0�U���U���E����u�U��U�E���$�p�M��U���U�M��Q�4�}  %�  �� +E�UԉE��U�}� |�}� r�U�+�E���E�"�M�-�U���U�E��؋M�� �ىE��M�U�U��E�� 0�}� |M	�}��  rBj h�  �M�Q�U�R�+|  ����0�M��U���Uj h�  �E�P�M�Q�C{  �E��U�U;U�u�}� |D�}�dr<j jd�E�P�M�Q��{  �Ѓ�0�E��M���Mj jd�U�R�E�P��z  �E��U�M;M�u�}� |D�}�
r<j j
�U�R�E�P�{  �ȃ�0�U�
�E���Ej j
�M�Q�U�R�z  �E��U��E���0�M��U���U�E�  �E�    �M�������E���]��������̋�U��EP�MQ��{  ��]���������̋�U���D�t�3ŉE��E�E܍M̉M��E�    j�U�R�E�P�M܋QR�P�t  ��3Ƀ} ���Mă}� u!h =j h*  h�<j�6  ����u̃}� u3�!Z  �    j h*  h�<h�>h =�B  ���   ��   3�;E��ىM�u!hx<j h+  h�<j�M6  ����u̃}� u3�Y  �    j h+  h�<h�>hx<�HB  ���   �   �}�u�E�E���M�3҃9-�E+E��M�Q�U��EBP�M�Q�U�3��:-��EP�p  ���Eȃ}� t�M� �E��$�URj �E�P�MQ�UR�EP�"   ���EȋEȋM�3�������]�����������̋�U���4�E�H���M��UR�M�� ���3��} ���E�}� u!h =j h�  h�<j�&5  ����u̃}� u@�X  �    j h�  h�<h�>h =�!A  ���E�   �M��o����E��  3�;U��؉E�u!hx<j h�  h�<j�4  ����u̃}� u@�X  �    j h�  h�<h�>hx<�@  ���E�   �M�������E��B  �U��t7�E3Ƀ8-��M�M��U�;Uu�E�E��E܋M��0�U܃��U܋E��  �M�M��U�:-u�E�� -�M����M��U�z j�E�P�  ���M��0�U����U���E�M�H�M��} ��   j�U�R��  ���M��r���� ���   ��E��
��U����U��E�x }]�M��t�U�B�؉E�&�M�Q��9U}�E�E���M�Q�ډŰẺE�MQ�U�R�W  ���EPj0�M�Q�ŝ�����E�    �M������EЋ�]������������̋�U���P�t�3ŉE��E�    �E�E��E� �MȉM�j�U�R�E�P�MċQR�P�np  ��3Ƀ} ���M��}� u!h =j ho  h�<j�2  ����u̃}� u3�V  �    j ho  h�<h?h =�>  ���   �i  3�;E��ىM�u!hx<j hp  h�<j�92  ����u̃}� u3�U  �    j hp  h�<h?hx<�4>  ���   �  �E؋H���M܋U�3��:-��E�E��}�u�M�M���U�3��:-���M+ȉM��U�R�EP�M�Q�U�R�l  ���E��}� t�E�  �E��   �M؋Q��9U����E��M؋Q���U܃}��|�E�;E|&�MQj�U�R�EP�MQ�UR�EP�_������D�B�M���t�U���M����M���t��U��B� �EPj�M�Q�UR�EP�MQ�������M�3�茙����]��������̋�U��Q�E�    �}et�}Eu%�E P�MQ�UR�EP�MQ�UR�
������E��{�}fu!�E P�MQ�UR�EP�MQ�c������E��T�}at�}Au%�U R�EP�MQ�UR�EP�MQ�2������E��#�U R�EP�MQ�UR�EP�MQ�������E��E���]Ë�U��j �EP�MQ�UR�EP�MQ�UR������]�������̋�U��} t#�EP�,:  ����P�MQ�UUR�uo  ��]Ë�U��Q�E�    �	�E����E��}�
s�M��� �R� �M��� ��ԋ�]���������������������������������̋�U���(  �������������5���=��f���f���f���f���f�%��f�-�������E ����E����E����������(�  ���������	 ����   �t��������x�������� � �j��R  ��j �� h$?�� �= � u
j�R  ��h	 ��� P�� ��]��̋�U���`�t�3ŉE��E� �E� �E� �E� �E� �E� �E���E��E���E���E���E���E���E���E���E��E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E� �E���E���E���E���E���E���E���E���E���E���E� �E� �E� �E� �E� �E� �E� �E׀�=�� t���P� �E���E�p�M��M؋U�U��}��  4�}��  ��  �E����E��}��   ��  �M���8� �$��� �E�-�  �E��}���  �M��$�� �E�   �E��@�U��]��E� �]��M��]ȍU�R�U؃���u�<P  � "   �E�E���c  �E�   �E��@�M��]��U��]��E� �]ȍM�Q�U؃���u��O  � !   �U�E���  �E�   �E��@�E� �]��M��]��U��]ȍE�P�U؃���u�O  � "   �M�E����  �E�   �E��@�U��]��E� �]��M��]ȍU�R�U؃���u�XO  � !   �E�E���  �E�   �E��@�M��]��U��]��E� �]ȍM�Q�U؃���u�O  � "   �U�E���3  �E�   �E��@�E� �]��M��]��U��]ȍE�P�U؃��M�E����  �E�   �E��@�U�����  �E�   �E��@�E� �]��M��]��U��]ȍE�P�U؃���u�iN  � "   �M�E���  �E�   �E��@�U��]��E� �]��M��]ȍU�R�U؃��E�E���S  �E�   �E��@�M��]��U��]��E� �]ȍM�Q�U؃���u��M  � "   �U�E���  �E�   �E��@�E� �]��M��]��U��]ȍE�P�U؃���u�M  � !   �M�E���  �E�   �E��@�U��]��E� �]��M��x"�U��E� �]��M��]��U��]ȍE�P�U؃���u�(M  � !   �M�E���O  �E�   �E��@�U��]��E� �]��M��]ȍU�R�U؃���u��L  � !   �E�E���  �E�   �E��@�M��]��U��]��E� �]ȍM�Q�U؃���u�L  � !   �U�E���  �E�   �E��@�E� �]��M��]��U��]ȍE�P�U؃���u�DL  � "   �M�E���k  �E�   �E��@�U��x"�E��M��]��U��]��E� �]ȍM�Q�U؃���u��K  � !   �U�E���  �E�   �E��@�E� �x"�M��U��]��E� �]��M��]ȍU�R�U؃���u�K  � !   �E�E���  �E�   �E��@�M��x"�U��E� �]��M��]��U��]ȍE�P�U؃���u�0K  � !   �M�E���W  �E�   �E��@�U��x"�E��M��]��U��]��E� �]ȍM�Q�U؃���u��J  � !   �U�E����  �E�   �E��@�E� �x"�M��U��]��E� �]��M��]ȍU�R�U؃���u�xJ  � !   �E�E���  �E�   �E�|@�M��x"�U��E� �]��M��]��U��]ȍE�P�U؃���u�J  � !   �M�E���C  �E�   �E��@�U��]��E� �]��M��]ȍU�R�U؃���u��I  � !   �E�E����  �E�   �E�t@�M��x"�U��E� �]��M��]��U��]ȍE�P�U؃���u�tI  � !   �M�E���  �E�   �E��@�U��]��E� �]��M��]ȍU�R�U؃���u�(I  � !   �E�E���O  �E�   �E��@�M��]��U��]��E� �]ȍM�Q�U؃���u��H  � !   �U�E���  �E�   �E�p@�E� �M�M��U��]��E� �]��M��]ȍU�R�U؃���u�H  � !   �E�E���   �E�   �E�l@�M��M�U��E� �]��M��]��U��]ȍE�P�U؃���u�*H  � !   �M�E���T�E�   �E�h@�U��M�E��M��]��U��]��E� �]ȍM�Q�U؃���u��G  � !   �U�E���M�3��܌����]�;� �� Ӣ � k� �� � Z� �� �� � /� � �� 3� �  	
�I ۦ 7� �� � K� �� � O� �� � @� �� ��U��j
�� ���3�]����������̋�U���h��  �(�P�  ���E��M���  ���  ��   ���E�$�  ���E�}� ~C�}�~�}�t�5h��  �U�R�V  ���E��   �E�P���E�$j�  ���   �M�Q�E�x"���$���E�$jj��  ���}���E�$�j  ���]��E��E������Dzh��  �U�R��  ���E��D�B�E��� th��  �M�Q�  ���E��$�"�U�R���E��$���E�$jj�K  ����]����̋�U��j
�� ���3�]�����������f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U��������̋�U��=�� u0�EP���E�$�����$���E�$�MQj�	  ��$�!��D  � !   h��  �UR�I  ���E]�̋�S�܃������U�k�l$���   �t�3ŉE��C P�KQ�SR�'  ����u)�E�����E��KQ�SR�CP�KQ�S R�E�P��  ���KQ�.
  ����|����=�� u>��|��� t5�S R���C�$�����$���C�$�CP��|���Q�  ��$�%���|���R�B	  ��h��  �C P�a  ���C�M�3��1�����]��[����������̋�U����E�@    �M�A    �U�B    �E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U��t�E��  ��E�H���U�J�E��t�E��  ��M�Q���E�P�M��t�E��  ��U�B���M�A�U�������������M�Q���ЋE�P�M�����҃������E�H���ʋU�J�E�����Ƀ������U�B�����M�A�U�������������M�Q���ЋE�P�M��� ��҃����E�H���ʋU�J�
  �E��E���t�M�Q���E�P�M���t�U�B���M�A�U���t�E�H���U�J�E���t�M�Q���E�P�M��� t�U�B���M�A�U�%   �E�}�   w�}�   t+�}� tI�}�   t.�K�}�   t�@�M����E��1�M�������E���M�������E���M�����E��M���   �U�t5�}�   t�}�   t�1�E����U�
�"�E������U�
��E������U�
�E%�  ���M��� ��ЋE��}  tT�M�Q ���E�P �M�Q ���E�P �M�U��Y�E�H`���U�J`�E�H`���U�J`�E�M��XP�X�U�B ���M�A �U�B �����M�A �U�E� �Z�M�Q`���E�P`�M�Q`�����E�P`�M�U��YP�  �EPjj �M�Q� �U�B����t�M�����E��M�Q����t�E�����U�
�E�H����t�U�����M��U�B���t�M����E��M�Q��t�E���ߋU�
�E����M�}�wb�U��$�ȴ �E���������   �U�
�@�E���������   �U�
�(�E���������   �U�
��E��������U�
�E������M�t�}�t�}�t.�;�U�%����   �M��%�U�%����   �M���U�%�����M��}  t�U�E�@P���M�U�BP���]�=� %� � �� �������̋�U��j �EP�MQ�UR�EP�MQ�UR������]�������̋�U���D�E���E��M��t �U��tj��  ���E�����E��  �M��t �U��tj��  ���E�����E��s  �M���   �U���  j�  ���E%   �E��}�   w�}�   tW�}� t �}�   tv��   �}�   ��   �   �M�������z���]�������]؋U�E���   �E�������z���]���(����]ЋM�E���Z�U�������z�(��]�������]ȋE�E���,�M�������z�(��]���(����]��U�E���E�����E��G  �M���;  �U���/  �E�    �E��t�E�   �M���������D��   �U�R�E��� �$�  ���]�M��   �M��}�����}�E��p"�]��E�   �   ���]�����Au	�E�   ��E�    �U��U��E��f�E��M��f�M��	�U����U��}����}:�E��t�}� u�E�   �M���M�U��t�E�   ��E�M���M�봃}� t�E����]�U�E����E�   �}� t
j�H  ���E�����E��M��t�U�� tj �%  ���E����E�3��}� ����]������������̋�U��� �EP��   ���E�}� t^�M�M��U�U�E�E�M�M��U�U�E �E��M$�M�h��  �U(R�{  ���E�P��^  ����u�MQ�/   ���E��"� h��  �U(R�G  ���EP�   ���E ��]�̋�U��Q�E�E��}�t�}�~ �}�~���9  � !   ��9  � "   ��]����̋�U��Q�E�    �	�E����E��}�}�M���0�;Uu�E���4����3���]���������������̋�U��Q�E�� t	�E�   �K�M��t	�E�   �:�U��t	�E�   �)�E��t	�E�   ��M��t	�E�   ��E�    �E���]�������̋�U����E�]��E�  �E��M���  �U����f�M��E���]����������̋�U��}  �u�} u�   �X�}  ��u�} u�   �B�E%�  =�  u�   �+�M���  ���  u�U����u�} t�   �3�]�����������̋�U����E��������Dz���]��E�    ��   �E%�  ��   �M����u
�} ��   �E�������]����Au	�E�   ��E�    �U�U��E��u/�M��M�U��   �t	�E���E�M��M�U����U����E%��  f�E�}� t�M�� �  f�Mj ���E�$�d������]��.j ���E�$�L������]��U���  ����-�  �E��M�U���E���]���������������̋�U��Q��}��E���]��������������̋�U��Q�}����E���]�������������̋�U�����}��E#E�M��U��#��f�E��m��E���]��̋�U����E��t
�-@��]���M��t����-@��]������U��t
�-L��]���E��t	�������؛�M�� t���]����]���������̋�U��j�hX�h � d�    P���SVW�t�1E�3�P�E�d�    �e�=�� ��   �E��@tp�=X� tg�E�    �U�E������Q�M���E�}�  �t�}�  �t	�E�    ��E�   �E�Ëe��X�    �M�ΈM�U�E�������U�⿉U�U�M�d�    Y_^[��]��������U���0���S�ٽ\�����=�� t��  ��8����   [����ݕz������U���U���0���S�ٽ\����=�� t�#  ��8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8����3  �   [�À�8�����=<� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �XA�����������HA����s4�hA�,ǅr���   �PA�����������@A����v�`AVW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�3X  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�����K   ����[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[��������̀zuf��\���������?�f�?f��^���٭^�����A�剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�����A�剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp�����A���۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-pA��p��� ƅp���
��
�t��������̋�U��Q�E�    �`���t
j
��   ���:A  �E��}� t
j�=  ���`���tjh  @j��  ��j�$�����]Ë�U��j�$W  ����tj�W  ����u#�=8�uh�   �k   ��h�   �^   ��]���������̋�U��Q�E�    �	�E����E��}�s�M��U;� Ju�E���$J���3���]���������������̋�U���   �t�3ŉE�EP�������E��}� ��  �E�    �}�   tN�}�   tE�}t?�M�Qj j j j�  �������������� t������t���E�   ��E�   �}� ��  j��U  ����tj��U  ������   �=8���   j��\ �E�}� tq�}��tk�E�    �	�U���U�}��  s%�E�M�U��J�������U�E��P��u����E� j �U�R������P�  ��P������Q�U�R�� ��  �}�   ��  ǅ����2�������- ����  +ȉ�����������������j h  hXNh@Nh�Mh\Mh  h ���_  ��P������3�������f��  h  ������Rj �� ��u:j h  hXNh@Nh�Lh�L������P������Q�_  ��P�t����������R�E_  ������<vk������P�._  ���������TA�������j h  hXNh@Nh8Ljh0L������+�������������+�Q������R��Z  ��P��~����j h  hXNh@Nh�Kh�Kh  h ��V  ��P�~����j h  hXNh@Nh K�E�Ph  h ��pV  ��P�~����h  h�Jh ��0T  ���M�3���q����]���������������̋�U��E�(�]�̋�U��E�U��DV�u�     j�E�P3�NVf�
�� ��u3�^��]ËM�U�E�QRP�� ��t�U��MZ  f9
u֋B<��~�8PE  u��HSW�x�D$+�3�3ۅ�t�;�r	��+�;p�rC��(;�r�;�t[C�=0� u �=,� uH�  �,���t:�0���,�h�NP�  3�;�t�U�R�UVV�M�QVVVR�Ѓ� ��u	_[3�^��]ËM����u���=��1��  �M���@�U�Rh�NV�Ѕ��p  �M��R VVV�E�PWS�҅��K  �M�u���@h�U�R�Є��(  �M�;��  ��B�Ѕ���   �M���Rj �E�P�E�P�EP�E�Pj �҄���   �E;�u�E�;�wE�;�r�M���B�Ѕ�u��   �E�����   =�����   ��    Qj �� P�� �����   �M���RV�E�Pj j j �E�P�҄�tR+}�;>rK�M��   ;�v
;<�r@;�r��D���Mj %��� ��M��Rpj j �EP�EP�E�P�҄�t�E�   Vj �� P�� �M����ҋM��P@�ҋM��P8�ҋM���P(�ҋE�_[^��]��������̋�U���  �t�3ŉE��=1� t3��M�3���n����]�V�5$ h�N�1��օ���  h�O�֋���u^�M�3��n����]�W�=  h�OV�׉�������u_^�M�3��tn����]�Sh�OV�׋؅�t4h|OV�׋���t&������Pjj h Oh  ���������tV�� [_3�^�M�3��n����]Í�����Q������������R������Pj h�NQǅ����  �Ӌ�����R����V�� ��u�������u��������u����r�Hf9�E����u�f��E����\t�\   f��E����@���+Ѓ��\����H��  �M�����N��N��E�������N�H��N�P��N�H��N�Pf��N�Hf�P������P�$ [_�M�3�^�m����]�����̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�   ���E��E�    �E���]�̋�U��EP�MQ�UR�EP�MQ�UR��\  ��]���������̋�U��P  ��q  �t�3ŉE��E�    �E�    �} u
�   �  ƅ���� h  ������Pj �p ��u8j h<  h Ph�Sh@Sh(Sh  ������Q��
  ��P�x�����������U��E�P�  ����@v]�M�Q�  ���U��D��E�j hE  h Ph�ShHRj�d�Q�U�������+й  +�Q�U�R�Go  ��P�x�����} t'�EP�<  ����@v�MQ�+  ���U�DÉE��I&  ��������<&  �     �}uǅ�����Q�
ǅ���� )�U���t�M�������
ǅ���� )�U���t�}uǅ�����Q�
ǅ���� )�M���tǅ�����Q�
ǅ���� )�} t�E�������
ǅ���� )�} tǅ�����Q�
ǅ���� )�} t�M�������
ǅ���� )�} tǅ�����Q�
ǅ���� )�}� t�U��������'�} t�E�������
ǅ���� )�������������}� tǅ�����O�
ǅ���� )�} tǅ�����Q�
ǅ���� )������R������P������Q������R������P������Q������R������P������Q������R������P�M�Q�U���OPhHQh�  h   ������Q� (  ��D�E�}� }*j h`  h Ph�Sh�8j"j�5$  �R�-����� �%$  ��������}� }8j he  h Ph�Sh�Ph�Ph   ������R��  ��P�u����h  h`P������P�ij  ��������������uj�0  ��j�6���������u�   �3��M�3��h����]������̋�U����E�E��M�Q�UR�EP�MQ�UR�EP�   ���E��E�    �E���]�̋�U��EP�MQ�UR�EP�MQ�UR�`  ��]���������̋�U��X"  �Qm  �t�3ŉE��E�    �E�    �} u
�   �  3�f������h  ������Qj �� ��u8j h<  h Ph�Wh@Wh�Lh  ������R�<T  ��P�#t�����������E��M�Q��S  ����@v`�U�R��S  ���M��TA��U�j hE  h Ph�WhHRj�h�P�M�������+����  +���P�M�Q��j  ��P�s�����} t'�UR�wS  ����@v�EP�fS  ���M�TA��U���!  � ��������!  �     �}uǅ����XV�
ǅ����TV�M���t�E�������
ǅ����TV�M���t�}uǅ����8V�
ǅ����TV�E���tǅ�����K�
ǅ����TV�} t�U�������
ǅ����TV�} tǅ����(V�
ǅ����TV�} t�E�������
ǅ����TV�} tǅ����V�
ǅ����TV�}� t�M��������'�} t�U�������
ǅ����TV�������������}� tǅ����0L�
ǅ����TV�} tǅ����V�
ǅ����TV������Q������R������P������Q������R������P������Q������R������P������Q������R�E�P�M��TRhXUh�  h   ������P�kj  ��D�E�}� }*j h`  h Ph�Wh�8j"j��  �Q踛���� �  ��������}� }8j hc  h Ph�Wh�ThhTh   ������P�&Q  ��P�q����h  h T������Q�F  ��������������uj�;,  ��j�����������u�   �3��M�3��5d����]�̋�U����E�    �E�    �	�E����E��}�$}Z�M��<�t�uK�U�k���8��E���p��M����M�h�  �U���p�P�` ��u�M���p�    3��뗸   ��]������̋�U����E�    �	�E����E��}�$}O�M��<�p� t@�U��<�t�t3�E���p��M��U�R�l j�E�P�T������M���p�    ��E�    �	�U����U��}�$}3�E��<�p� t$�M��<�t�u�U���p��E�M�Q�l 뾋�]��̋�U��j�hx�h � d�    P���SVW�t�1E�3�P�E�d�    �E�   �=�� u�����j������h�   �������E�<�p� t
�   �   h  h�Wjj�w�����E�}� u�'  �    3��   j
�   ���E�    �M�<�p� uDh�  �U�R�` ��u"j�E�P��������  �    �E�    ��M�U��p��j�E�P�݂�����E������   �j
�e   ��ËE��M�d�    Y_^[��]������������̋�U��E�<�p� u�MQ��������u
j�������U��p�P�� ]�̋�U��E��p�Q�� ]��������̋�U���(�} t�} v	�E�   ��E�    �E�E�}� uhYj jh�Xj�K�������u̃}� u0�  �    j jh�Xh�XhY�I  ���   �L  �} ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U�E�Ph�   �M��Q�@b����3҃} �U��}� uhdXj jh�Xj��������u̃}� u0��  �    j jh�Xh�XhdX�  ���   �  �M�M��U�U��E��M���E���U����U��E���E��t�M����M�t�̓}� ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�<a�����<X��t3�t	�E�   ��E�    �M܉M�}� uh Xj jh�Xj�k�������u̃}� u-��  � "   j jh�Xh�Xh X�i  ���"   �o�}�tg�}���t^�E+E���;EsP�M+M����U+�9��s
����E���M+M����U+щU؋E�Ph�   �M+M��U�D
P�U`����3���]������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+������̋�U��Q�E�    �}�wC�EP�t   ���E��}� t�*�=�� u�h  �    ��MQ��  ����u����UR�  ���9  �    3���}� u�$  �    �E���]�������̋�U��Q�=�� u�l���j������h�   �h������} t�E�E���E�   �M�Qj ���R�� ��]���������̋�U��QV�E�    �} u�4�EPj ���Q�� �E��}� u�D P��  �����h  �0^��]�̋�U��E���]�̋�U��Q����E��M�Q� �E��}� t�UR�EP�MQ�UR�EP�U�����MQ�UR�EP�MQ�UR�
   ��]������̋�U��jh �j�   ��h ��� P�� ]������̋�U���8  �t�3ŉE��}�t�EP�\  ��ǅ����    jLj ������Q�]�����������U��� ����E��E�    ǅ���    ������������������������������������f������f������f������f������f������f�������������ǅ ���  �M�������U�������E�H��������U�������E�������M������� �E�j �� �U�R�� ���������� u�}� u�}�t�EP�B  ���M�3��Z����]��SVW�T$�D$�L$URPQQh�� d�5    �t�3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�Bf  �   �C�Tf  �d�    ��_^[ËL$�A   �   t3�D$�H3���Y��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�e  3�3�3�3�3���U��SVWj Rhv� Q��6 _^[]�U�l$RQ�t$������]� �������������̋�U��Q�EP�< �M���    t�U���   P�< �M���    t�U���   P�< �M���    t�U���   P�< �M���    t�U���   P�< �E�    �	�M����M��}�m�U����E�|H��t$�M����U�|
P t�E����M�TPR�< �E����M�|L t$�U����E�|T t�M����U�D
TP�< 넋M���   �´   R�< ��]�̋�U��Q�} �  �EP�H �M���    t�U���   P�H �M���    t�U���   P�H �M���    t�U���   P�H �M���    t�U���   P�H �E�    �	�M����M��}�m�U����E�|H��t$�M����U�|
P t�E����M�TPR�H �E����M�|L t$�U����E�|T t�M����U�D
TP�H 넋M���   �´   R�H �E��]����̋�U��Q�E���    ��   �M���   ȼ��   �U���    ��   �E���   �9 ��   �U���    t4�E���   �9 u&j�U���   P�zw�����M���   R��i  ���E���    t4�M���   �: u&j�E���   Q�:w�����U���   P��h  ��j�M���   R�w����j�E���   Q� w�����U���    to�E���   �9 uaj�U���   -�   P��v����j�M���   ��   R�v����j�E���   ��   Q�v����j�U���   P�v�����M���   ��t8�U���   ���    u&�M���   R�a  ��j�E���   Q�>v�����E�    �	�U����U��}���   �E����M�|H��t:�U����E�|P t*�M����U�D
P�8 uj�M����U�D
PP��u�����M����U�|
L t�E����M�|T uA�U����E�|L u�M����U�|
T t!h�`j h�   h�`j���������u̋M����U�|
L t:�E����M�|T t*�U����E�LT�9 uj�U����E�LTQ�*u���������j�UR�u������]Ë�U��Q�} t�} u3��\�E��M��U�;UtI�E�M��UR�������}� t�E�P�������}� t�M��9 u�}� �t�U�R�������E��]����������̋�U��j�h��h � d�    P���SVW�t�1E�3�P�E�d�    �Ie���E��E��Hp#t�t	�U��zl uDj�������E�    �صP�M���lQ�������E��E������   �j����������d���Pl�U�}� u
j 胋�����E�M�d�    Y_^[��]�����������̋�U��j�h��h � d�    P���SVW�t�1E�3�P�E�d�    �yd���E��E��Hp#t�t�U��zl ��   j��������E�    �E��Hh�M�U�;�tI�}� t%�E�P�H ��u�}��tj�M�Q�s�����U���Bh���M�U�R�< �E������   �j��������	�E��Hh�M�}� u
j �l������E�M�d�    Y_^[��]����̋�U��j�hؠh � d�    P���SVW�t�1E�3�P�E�d�    �E������bc���E������E܋Hh�M��UR�H  ���E�E��M;H�  hN  h�ejh   ��e�����E��}� ��  �U܋rh��   �}��E��     �M�Q�UR��  ���E؃}� ��  �E܋HhQ�H ��u�U܁zh�tj�E܋HhQ�q�����U܋E��Bh�M܋QhR�< �E܋Hp���-  �t����  j��������E�    �E��H����U��B����M��Q����E�    �	�E���E�}�}�M�U�E�f�TPf�M�����E�    �	�E���E�}�  }�M�M�U�A�� ����E�    �	�M���M�}�   }�U�U�E䊊  ����׋�R�H ��u�=��tj��P�p�����M����U�R�< �E������   �j��������(�}��u"�}��tj�E�P�Kp�����
  �    ��E�    �E؋M�d�    Y_^[��]���������������̋�U��j�hhd�    P��$�t�3�P�E�d�    �E�    �E�P�M������E�    ���    �}�u)���   �� �E��E������M��}����E��}�c�}�u)���   �� �E��E������M��N����E��N�4�}�u.���   �M��_�����Q�U��E������M������E���E�E��E������M������EЋM�d�    Y��]������������̋�U���,�t�3ŉE�V�EP��������E�} u�MQ�  ��3���  �E�    �	�U����U��}��E  �E�k�0���;M�+  �E�    �	�U����U��}�  s�EE��@ ���E�    �	�M����M��}�s{�U�k�0�E���� ��M��	�U���U�E����tN�U��B��tC�M���U��	�E����E��M��Q9U�w!�E�����UU��B��MM��A����v����U�E�B�M�A   �U�BP�  ���M�A�E�    �	�U����U��}�s�E�k�0�M��U�u�f��p�f�DJ�ӋMQ�#  ��3��  �����} t!�}��  t�}��  t�UR�� ��u����k  �E�P�MQ�� ���9  �E�    �	�U����U��}�  s�EE��@ ��M�U�Q�E�@    �}���   �MމM��	�Uԃ��UԋE����tE�U��B��t:�M���U��	�E����E��M��Q9U�w�EE��H���UU��J����E�   �	�E����E��}��   s�MM��Q���EE��P�֋M�QR�   ���M�A�U�B   �
�E�@    �E�    �	�M����M��}�s3ҋE��Mf�TA��UR�  ��3���=�� t�EP�   ��3�����^�M�3��J����]�����������̋�U��Q�E�E��M���  �M��}�w-�U����� �$��� �  ��  ��  �	�  �3���]ÍI _� f� m� t� {�  ����̋�U��Q�E�    �	�E����E��}�  }�MM��A ��U�B    �E�@    �M�A    �E�    �	�U����U��}�}3��M��Uf�DJ���E�    �	�E����E��}�  }�MM��U������A���E�    �	�M����M��}�   }�UU��E�������  �׋�]���������̋�U���(  �t�3ŉE�������P�M�QR�� ���-  ǅ����    ���������������������   s��������������������ƅ���� ������������������������������������tD�����������������������������������Q9�����w������Ƅ���� ���j �M�QR�E�HQ������Rh   ������Pjj �`  �� j �M�QRh   ������Ph   ������Qh   �U�BPj �]  ��$j �M�QRh   ������Ph   ������Qh   �U�BPj ��\  ��$ǅ����    ���������������������   ��   ��������U������t:�M������Q���E������P�M�������������������  �]��������M������t:�E������H�� �U������J�E�������������������  ��E�����ƀ   �2�����   ǅ����    ���������������������   ��   ������Ar?������Zw6�U������B���M������A�������� �E�������  �X������ar?������zw6�M������Q�� �E������P�������� �U�������  ��E�����ƀ   �<����M�3��F����]����̋�U��=�� uj��K��������   3�]����������̋�U��V��   �M��UR�   �����   �0^]��������̋�U��Q�E�    �	�E����E��}�-s�M��U;� �u�E�����7�ԃ}r�}$w	�   �"� �}�   r�}�   w	�   ���   ��]������������̋�U��Q�UV���E��}� u	�h����E�����]���������̋�U��Q�%V���E��}� u	�l����E�����]���������̋�U��E���]�̋�U��Q���P� �E��}� t�MQ�U�����u3���   ��]����������̋�U��   ]����̋�U�����    ]���������������̋�U���V3��} ���E�}� uh�fj jHh0fj�p�������u̃}� u-������    j jHh0fhfh�f�n�����3��   �}�v�����    3��~�} u�E   �URj ���P�� �E��MQ�URj���P�� �E��}� u:�}� @  w�M;M�w�8   ��t�U�U���D P���������&����0�E�^��]������������̋�U����E�����j j�E�Pj ���Q�� ��t�}�u	�E�   ��E�    �E���]���������̋�U���V�E�E��} u�MQ��������   �} u�UR�������3��   �E�    �}�w)�} u�E   �EP�MQj ���R�� �E���EP�������:����    3��e�}� u	�=�� u%�}� t��D P�������������0�E��1�MQ�c�������u�D P�`�������������03���J���^��]������̋�U��Q�E�����j j ���P�L ��u�E������E���]�̋�U��Q�E�E��M�Qj �UR�EP�MQ�M]  ����]������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�_  ����]��̋�U��E��=   vhgj j8h�fj��������u̋UR�EPj �   ��]������������̋�U����EP�M���q���M����   vhgj jDh�fj�)�������u̃}�|5�}�   ,�M���r��� ���   �U�Q#E�E�M��|r���E��1�'�M��r������   �B�#E�E�M��Sr���E���M��Fr����]��̋�U���(�EP�M��Lq���}�|6�}�   -�M��Er������   �E�B#M�M��M���q���E��   �M��r��P�U�����   R��a  ����t!�E��%�   �E�M�M��E� �E�   ��U�U��E� �E�   j�M���q��� �HQ�M��q����BP�M�Q�U�R�E�Pj�M��q��P��W  �� ��u�E�    �M��Lq���E���M�#M�M؍M��5q���E؋�]���������������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u��a  ��   u������r)��$�� �Ǻ   ��r����$�$� �$� � ��$��� �4� `� �� #ъ��F�G�F���G������r���$�� �I #ъ��F���G������r���$�� �#ъ���������r���$�� �I � �� �� �� �� �� �� �� �D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�� �� � (� 4� H� �E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��� �����$�\� �I �Ǻ   ��r��+��$��� �$��� ��� �� � �F#шG��������r�����$��� �I �F#шG�F���G������r�����$��� ��F#шG�F�G�F���G�������V�������$��� �I `� h� p� x� �� �� �� �� �D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��� ���� �� �� �� �E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_����������������̋�U����E�E��M����MZ  t3��;�E��M�H<�M�U�:PE  t3�� �E���E��M����  t3���   ��]�̋�U����E�MH<�M��E�    �U��B�M��T�U���E����E��M��(�M�U��B9E�s#�M�U;Qr�E�H�U�J9Ms�E���3���]�����������̋�U��j�h �h � d�    P���SVW�t�1E�3�P�E�d�    �e��E�   �E�    �E�P���������u�E�    �E������E��   �M+M�M܋U�R�E�P�������E��}� u�E�    �E������E��b�M��Q$��   ���҃��U��E������E��@�E������7�E���U؋E�3�=  �����Ëe��E�    �E������E���E������M�d�    Y_^[��]��������������̋�U��h0� � � �]���������̋�U��j�h@�h � d�    P���SVW�t�1E�3�P�E�d�    �e��fK���@x�E�}� t#�E�    �U��E�������   Ëe��E������"����M�d�    Y_^[��]Ë�U��Q�K���@|�E��}� t�U��a�����]�������������̋�U��j�h`�h � d�    P���SVW�t�1E�3�P�E�d�    �e� �P� �E�}� t#�E�    �U��E�������   Ëe��E�����������M�d�    Y_^[��]������������̋�U��E���M���U���E��]�����������������������̋�U��j�h��h � d�    P���SVW�t�1E�3�P�E�d�    �E�    �E�    �E�EċMă��Mă}���   �U�����$���E���MЋ�U�E؃��E��  �E���MЋ�U�E؃��E���   �E���MЋ�U�E؃��E���   �E���MЋ�U�E؃��E��   �}H���E��}� u�����  �M��Q\R�EP�  �����EЋMЋ�U��   �x3�t	�E�   ��E�    �M��Mȃ}� u!h�gj h�  hHgj�,�������u̃}� u1�����    j h�  hHgh�gh�g�'���������4  �E�P� �E�}�u3��  �}� uj��n���}� t
j ��������E�    �}t�}t�}u,�M��Q`�U܋E��@`    �}u�M��Qd�ŰE��@d�   �}u<�p;�M��	�Uԃ��Uԡp;t;9E�}�M�k��U��B\�D    ���
�	C���MЉ�E������   ��}� t
j �Y�����Ã}u�U��BdPj�U���
�MQ�U���}t�}t�}u�U��E܉B`�}u	�M��ỦQd3��M�d�    Y_^[��]Ë� � T q 7 �  ������̋�U��Q�E�E��M��Q;Ut�E����E��|;k�M9M�s�ً|;k�U9U�s�E��H;Mu�E���3���]����̋�U���P� ]�������������̋�U��E��]�̋�U��jj �EPj �   ��]�������̋�U��j�h�d�    P���t�3�P�E�d�    �EP�M��=e���E�    �M�M�M��7f���P�E�L#Mu;�} t�M��f������   �M�H#U�U���E�    �}� u	�E�    ��E�   �E؉E��E������M��e���E��M�d�    Y��]��������������̋�U����E%�����E�M#M��������   �} tj j �|W  ���U�3�t	�E�   ��E�    �M��M��}� uh�hj j1hhj��������u̃}� u-������    j j1hhh�gh�h�}������   �/�} t�EP�MQ��V  ���U���EP�MQ��V  ��3���]Ë�U����EP�M��c���M��d����t/�M��d������   ~�M��d��Pj�UR�������E��j�EP�M��sd��P�M������E�M�M�M��)d���E��]��̋�U��=P� uj�EP���������j �MQ�U�����]Ë�U���4�EP�M���b���}   ��   �M���c����t/�M���c������   ~�M���c��Pj�UR�\������E��j�EP�M��c��P�������Ẽ}� t,�M��c������   �E��M��M��Rc���E��*  ��U�U܍M��:c���E��  �M��Zc��� ���   ~D�M��Gc��P�M�����   Q�S  ����t"�U�����   �U��E�E��E� �E�   ������� *   �M�M��E� �E�   j�M���b����BPj�M�Q�U�R�E�Ph   �M���b����QR�M��b��P�E  ��$�E�}� u�E�E؍M��fb���E��A�}�u�M��MԍM��Lb���E��'��U��E���ЉUЍM��-b���E���M�� b����]������������̋�U��Q�=P� u$�}A|�}Z�E�� �E���M�M��E���j �UR���������]�����������̋�U���@�t�3ŉE��E�    �E�    �EP�M��`���M��a��Pj j j j �MQ�U�R�E�P��`  �� �E��MQ�U�R�Z  ���E��E���u8�}�u�E�   �M��<a���E��j��}�u�E�   �M�� a���E��N�:�M���t�E�   �M��a���E��0��U���t�E�   �M���`���E���E�    �M���`���E��M�3���.����]���������������̋�U���@�t�3ŉE��E�    �E�    �EP�M��_���M��`��Pj j j j �MQ�U�R�E�P��_  �� �E��MQ�U�R�_  ���E��E���u8�}�u�E�   �M��,`���E��j��}�u�E�   �M��`���E��N�:�M���t�E�   �M���_���E��0��U���t�E�   �M���_���E���E�    �M���_���E��M�3���-����]���������������̋�U����E�E��M�Q�U�3��} ���E�}� uh =j j7h`ij���������u̃}� u0�>����    j j7h`ihLih =��������   �$  3�;U��؉E�uhx<j j8h`ij�p�������u̃}� u0������    j j8h`ihLihx<�n������   ��  �U� 3��} ����#E��;E��ىM�uh�hj j=h`ij���������u̃}� u0�d���� "   j j=h`ihLih�h��������"   �J  3��} ���E�}� uh�hj j>h`ij��������u̃}� u0������    j j>h`ihLih�h�������   ��   �U��0�E����E��} ~A�M����t�E���M�U����U���E�0   �E��M��U����U��E���E빋M�� �} |>�U����5|3�M����M��U����9u�M��0�U����U���E�����U��
�E���1u�U�B���M�A�&�U��R���������P�E��P�MQ�$  ��3���]�����������̋�U���,�t�3ŉE��EP�M�Q�   ���U�Rj j���ċMԉ�U؉Pf�M�f�H�l  ���U�B�E�M��U��E�Pj j(h8jh$jh�i�M�Q�UR�EP�I�����P��6�����M�U�Q�E�M�3��W*����]���̋�U����E�   �3�f�E��M�Q���  ��f�U��E�H�� �  f�M�U�B%�� �E�M��U��E��E�}� t�}��  t�P��  f�M��a�}� u)�}� u#�U�B    �E�     �Mf�U�f�Q�   �E�<  f�E��E�    ��M����  f�M��U����?  f�U��E���E��M�����U�B�E����M��U�B%   �u;�M�Q��E���   ������ыE�P�M���E�f�M�f��f�M���U��E�ЋMf�Q��]��������������U��WV�u�M�}�����;�v;���  ���   r�=�� tWV����;�^_u�K  ��   u������r)��$�P�Ǻ   ��r����$�d�$�`��$���t��#ъ��F�G�F���G������r���$�P�I #ъ��F���G������r���$�P�#ъ���������r���$�P�I G4,$�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�P��`ht��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$���I �Ǻ   ��r��+��$���$��� $L�F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ���������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�����(�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�����������������SW3��D$�}G�T$���ڃ� �D$�T$�D$�}�T$���ڃ� �D$�T$�u�L$�D$3���D$���3�OyN�S�؋L$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$Oy���؃� _[� ��������������WVS3��D$�}G�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u�L$�D$3���؋D$����A�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�Ou���؃� [^_� �����̀�@s�� s����Ë�3������3�3��̀�@s�� s����Ë�3Ҁ����3�3���U��W�}3�������ك��E���8t3�����_����̋�U��j�D\����]���������������̋�U����} uh�kj jdh0kj轺������u̋M�M��U�R腀  ���E��E��H��   u$����� 	   �U��B�� �M��A����G  �-�U��B��@t"������ "   �M��Q�� �E��P����  �M��Q��tH�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J�����  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6�|  �� 9E�t�|  ��@9E�u�M�Q��{  ����u�U�R��z  ���E��H��  ��   �U��E��
+Hy!h�jj h�   h0kj�>�������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P� m  ���E��q�}��t!�}��t�M����U���������U���E����E��H�� t7jj j �U�R�oi  ���E�U�E�#E���u�M��Q�� �E��P����O�M��Q�E���E�   �M�Q�UR�E�P�bl  ���E�M�;M�t�U��B�� �M��A�����E%�   ��]����̋�U��E����U�
�E��A�]����̋�U��E����U�
�E��A��Q�]�̋�U��E����U�
�E�f�A�]���̋�U��3�]�������̋�U����E���]��E���]���������̋�S�܃������U�k�l$���   �t�3ŉE��C��M��U��U�C��M��U����U��}�w@�E��$�0�E�   �4�E�   �+�E�   �"�E�   ��E�   ��K�   �E�    �}� ��   �U�P�K��Q�U�R軜������ul�C�E�}�t�}�t�}�t� �M����M��U������U��C�@�]��	�M�����M��S��R�C��P�KQ�U�R�E�P��p���Q������h��  �U�P������ǅl���    �K�9t�=�� u�SR�q�������l�����l��� u�C�Q褟�����M�3������]��[��
�.%��U����E�    �E�E�}� |,�}�~�}�t��4��M��U�4��y�4��E��o3�t	�E�   ��E�    �U��U��}� uh�nj j9hpnj�d�������u̃}� u+������    j j9hpnhLnh�n�b����������E���]���̋�U���@�t�3ŉE��E�    ��*���E��E�    �E�    �E�    �= � ��   hlo�$ �Eԃ}� u3��  h`o�E�P�  �E��}� u3��  �M�Q� � �hPo�U�R�  P� �$�h<o�E�P�  P� �(�h o�M�Q�  �E��U�R� �0��=0� tho�E�P�  P� �,��,�;M�th�0�;U�t]�,�P� �EЋ0�Q� �Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W�$�;M�t�$�R� �Eȃ}� t�UȉE�}� t*�(�;E�t �(�Q� �Eă}� t
�U�R�UĉE� �P� �E��}� t�MQ�UR�EP�M�Q�U���3��M�3������]Ë�U���4�} t�} v	�E�   ��E�    �E�E�}� uh�pj jh(pj軲������u̃}� u0�'����    j jh(phph�p蹾�����   �\  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E��M���Qh�   �U��R�����3��} ���E��}� uhdXj jh(pj��������u̃}� u0�^����    j jh(phphdX�������   �  �U�U��E�E��}� v�M����t�E����E��M����M��܃}� ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E܋M���Qh�   �U��R�������o��t3�t	�E�   ��E�    �U؉U�}� uh�oj j h(pj��������u̃}� u0�N����    j j h(phph�o�������   �  �M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���MԋU���Rh�   �E��P������<X��t3�t	�E�   ��E�    �EЉE�}� uh Xj j*h(pj�ί������u̃}� u-�:���� "   j j*h(phph X�̻�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9��s����U���E+E����M+ȉM̋U���Rh�   �E+E��M�TAR�����3���]������������̋�U���,�} u�} u�} u3���  �} t�} v	�E�   ��E�    �E�E�}� uh�pj jh�pj貮������u̃}� u0�����    j jh�ph�ph�p谺�����   �`  �} u`3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E�M���Qh�   �U��R�����3���  �} ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P�>����3Ƀ} ���M��}� uhdXj jh�pj脭������u̃}� u0������    j jh�ph�phdX肹�����   �2  �E�E��M�M��}�u7�U��Ef�f�
�U���M����M��U���U��t�E����E�t���}�WM����t&�M;Mrh<Xj j+h�pj�֬������u̋E��Mf�f��E���U����U��E���E��t�M����M�t�U���Ut���} u3��M�f��}� ��   �}�u3ҋE�Mf�TA��P   �E  3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E܋M���Qh�   �U��R������<X��t3�t	�E�   ��E�    �U؉U�}� uh Xj j>h�pj���������u̃}� u-�-���� "   j j>h�ph�ph X迷�����"   �r�}�tj�}���ta�M+M���;MsS�U+U����E+�9��s����M���U+U����E+EԋM���Qh�   �U+U��E�LPQ�����3���]���������������̋�U��Q�E�E��M���E����E���t��E�+E������]Ë�U���(�} t�} v	�E�   ��E�    �E�E�}� uh�pj jh�Xj苪������u̃}� u0������    j jh�Xhdqh�p艶�����   �X  �} ��   3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E�M���Qh�   �U��R�|����3��} ���E��}� uhdXj jh�Xj�©������u̃}� u0�.����    j jh�XhdqhdX��������   �  �U�U��E�E��M��Uf�f��M���E����E��M���M��t�U����U�t�˃}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P�s�����<X��t3�t	�E�   ��E�    �E܉E�}� uh Xj jh�Xj袨������u̃}� u-����� "   j jh�Xhdqh X蠴�����"   �r�}�tj�}���ta�U+U���;UsS�E+E����M+�9��s����U���E+E����M+ȉM؋U���Rh�   �E+E��M�TAR�����3���]Ë�U��} t�E�M��U���U�E]���������������̋�U��Q�} tV�E���E�M��U��}���  u�EP�������.�}���  t%3�u!h�qj h�   hxqj�g�������u̋�]����������̋�U���]��������̋�U��j�hȡh � d�    P���PP  ��  �t�1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    ƅп�� h�  j ��ѿ��P�c����ƅ���� h�  j ������Q�F����3�f������h�  j ������P�'����ƅЯ�� h�  j ��ѯ��Q�
�����} |�}|����*  �E�    �}��   h���< ����   j h  h0rh�wh�wj
h   ��п��R�EP�z  ��P�)����hXw�� �} t�M�������
ǅ����Hw������R�� h@w�� ��п��P�� hT(�� �[���ǅ���������=  �} ��   ǅ̯��    �������ȯ��������     �UR�EPh�  h   ��Я��Q��/  ����̯����̯�� }*j h*  h0rh�wh�8j"j�����R�D���� ������ȯ�����̯�� }8j h-  h0rh�wh�vh�Ph   ��Я��R�D�����P�������}uV�} tǅ�����v�
ǅ����|vj h2  h0rh�wh�u������Ph   ��п��Q������P�����j h4  h0rh�whpu��Я��Rh   ��п��P��t  ��P�U�����}u�M������t8j h9  h0rh�wh(uh uh   ��п��P�t  ��P�����j h:  h0rh�wh�thT(h   ��п��Q�it  ��P�������} ��   ǅį��    ����������������     ��п��P�MQ�URh�th�  h   ������P�w�������į����į�� }*j hA  h0rh�wh�8j"j�����Q�B���� �������������į�� }8j hD  h0rh�wh�Ph�Ph   ������P�I�����P�������:j hH  h0rh�whpt��п��Qh   ������R������P�����ǅ����    ǅ����    j�������Ph   ������Q������R��r  ��������j hM  h0rh�wh�sj"j������P�A���� ������ t8j hO  h0rh�whsh�rh   ������Q�%�����P������=�� u�=�� �#  ǅ����    ǅ����    j�Ȩ�����E�   �����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   �������������렃����� un�����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���tǅ����   ���������������E�    �   �j������Ã����� �D  �=�� t?ǅ����    ������R������P�MQ�������tǅ����   ������������������ ��   �E������t>�U�<����t1j ������P������Q�m�����P������R�E����Q�� �U������t������Q�� �U������twƅп�� �} t9j h�  h0rh�wh�wj
h   ��п��Q�UR�,t  ��P�������Я��P�MQ�U��ҍ�п��#�R�MQ�UR�h������������E������   ��}uh���H Ë������M�d�    Y_^[�M�3�������]�������������̋�U��j�h�h � d�    P���\�  �  �t�1E�3ŉE�SVWP�E�d�    ǅ����    ǅ����    3�f��Я��h�  j ��ү��Q�1	����3�f������h�  j ������P�	����ƅ���� h�  j ������Q������3�f��Џ��h�  j ��ҏ��P�������} |�}|����.  �E�    �}��   h���< ����   j h�  h0rh�}h�}j
h   ��Я��Q�UR��  ��P������hP}�� �} t�E������
ǅ���0}�����Q�� h }�� ��Я��R�� h}�� �'���ǅ���������A  �} ��   ������ ��ȏ��������     �MQ�URh�  h   ��Џ��P�8�  ����̏����̏�� }*j h  h0rh�}h�8j"j�w����Q�o<���� �g�����ȏ�����̏�� }8j h  h0rh�}h�|hhTh   ��Џ��P�������P�������}uV�} tǅ���T|�
ǅ���0|j h  h0rh�}h�{�����Qh   ��Я��R�~�����P�e����j h  h0rh�}h {��Џ��Ph   ��Я��Q������P�+�����}u�U������t8j h  h0rh�}h�zh�zh   ��Я��Q�������P������j h  h0rh�}h�zh}h   ��Я��R������P������} ��   ǅď��    ����� �������ݾ���     ��Я��Q�UR�EPhhzh   h   ������Q�-	  ����ď����ď�� }*j h  h0rh�}h�8j"j�|����R�t:���� �l������������ď�� }8j h  h0rh�}h�ThhTh   ������R�������P�������:j h"  h0rh�}hz��Я��Ph   ������Q������P�����ǅ����    j h(  h0rh�}hxyj"jj�������Rh   ������Pj ��z  ��P�9���� ������������ t8j h*  h0rh�}h�xhtxh   ������Q�P�����P�������=�� u�=�� �#  ǅ����    ǅ����    j賠�����E�   �����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   �렃����� un�����������������H������������ tHǅ����    ������R������P�MQ�������B�Ѓ���t������������ǅ����   ���E�    �   �j������Ã����� �g  �=�� t?ǅ����    ������R������P�MQ�������t������������ǅ����   ������ �  �E�������[  �U�<�����J  �E����Q�d ����������t�Jj ������R������P�������P������Q�U����P�� ��t��   �D ��t��   ǅ���    j h{  h0rh�}h�wj"jj�������Qh   �����R�����P�4x  ��P��6���� ���������� t>�����Pt5j ������Q������R�+�������P������P�M����R�� �@����� v������������j ������Q�����R�����P�M����R�� �E������t������R�� �E������ty3�f��Я���} t9j h�  h0rh�}h�}j
h   ��Я��P�MQ�}  ��P�{������Џ��R�EP�M��ɍ�Я��#�Q�EP�MQ蠖�����������E������   ��}uh���H Ë������M�d�    Y_^[�M�3�������]�����̋�U���@�t�3ŉE��E�    ����E��E�    �E�    �E�    �=4� ��   hlo�$ �Eԃ}� u3��  h,~�E�P�  �E��}� u3��  �M�Q� �4�hPo�U�R�  P� �8�h<o�E�P�  P� �<�h~�M�Q�  �E��U�R� �D��=D� tho�E�P�  P� �@��@�;M�th�D�;U�t]�@�P� �EЋD�Q� �Ẽ}� t8�}� t2�UЉE�}� t�U�Rj�E�Pj�M�Q�U̅�t�U��u�E�   �}� t�E    �E�W�8�;M�t�8�R� �Eȃ}� t�UȉE�}� t*�<�;E�t �<�Q� �Eă}� t
�U�R�UĉE�4�P� �E��}� t�MQ�UR�EP�M�Q�U���3��M�3��d�����]Ë�U����} u3��k  3��} ���E��}� uh�~j j7h�~j脓������u̃}� u0�����    j j7h�~h|~h�~肟�����   �  �} t�U;U��   �EPj �MQ������3҃} �U��}� uhd~j j=h�~j���������u̃}� u-�f����    j j=h�~h|~hd~��������   �~�M;M҃��U�uh8~j j>h�~j虒������u̃}� u-����� "   j j>h�~h|~h8~藞�����"   ��   ��MQ�UR�EP赻����3���]�������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ������̋�U��Q�E�E��M�Qj �UR�EP�MQ�UR�9u  ����]���SV�D$�u�L$�D$3���؋D$����A�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$vN3ҋ�^[� ��������S�D$�u�L$�D$3���D$���3��P�ȋ\$�T$�D$���������u�����d$��d$�r;T$wr;D$v+D$T$+D$T$���؃� [� ����������̋�U��QS�E���E�d�    �d�    �E�]�m��c���[��]� ������������XY�$����������̋�U���SVWd�5    �u��E��>j �EP�M�Q�UR��  �E�H����U�Jd�=    �]��;d�    _^[��]� ������U���SVW��E�j j j �E�P�MQ�UR�EP�MQ�${  �� �E�_^[�E���]����̋�U����E�    �E�?�t��M�3��E��U�U�E�E��M���M�d�    �E�E�d�    �UR�EP�MQ腏  �E�E�d�    �E��]��̋�U��Q��E�H3M����j �MQ�U�BP�M�QRj �EP�M�QR�EP�az  �� �E��E���]����̋�U���8S�}#  u��@�M��   ��   �E�    �E��@�t��M�3��E��U�U�E�E�M�M�U �U��E�    �E�    �E�    �e�m�d�    �E؍E�d�    �E�   �E�E̋M�M��2	�����   �UԍE�P�M�R�Uԃ��E�    �}� td�    ��]؉d�    �	�E�d�    �E�[��]����̋�U��QS��E�H3M������M�Q��ft�E�@$   �   �v�tj�M�QR�E�HQ�U�BPj �MQ�U�BP�MQ��x  �� �U�z$ u�EP�MQ�6���j j j j j �U�Rh#  �~������E��]�c�k ��   [��]���̋�U��Q�} �E�HSV�pW�M�����|8����u�����E��MN��9L���};H~���u�M���ރ} }̋E�M�UF�1�:;xw;�v�м���M�_��^��[��]Ë�U��EV�u�������   �N������   ��^]����̋�U���v�����   ��t�M9t�@��u��   ]�3�]���̋�U��V�E���u;��   u�5���N���   ^]��$�����   �x t�H;�t���x u�^]�����V�P^]����������U��SVWUj j h�B�u�\�  ]_^[��]ËL$�A   �   t2�D$�H�3�����U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h Cd�5    �t�3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y Cu�Q�R9Qu�   �SQ����SQ����L$�K�C�kUQPXY]Y[� �����������̋�U��} u�W  j�E�HQ�����j�U�BP�����j�M�QR�����j�E�HQ�o����j�U�BP�^����j�M�QR�M����j�E�Q�=����j�U�B P�,����j�M�Q$R�����j�E�H(Q�
����j�U�B,P������j�M�Q0R������j�E�H4Q������j�U�BP������j�M�Q8R�����j�E�H<Q�����j�U�B@P�����j�M�QDR�����j�E�HHQ�q����j�U�BLP�`����j�M�QPR�O����j�E�HTQ�>����j�U�BXP�-����j�M�Q\R�����j�E�H`Q�����j�U�BdP������j�M�QhR������j�E�HlQ������j�U�BpP������j�M�QtR�����j�E�HxQ�����j�U�B|P�����j�M���   R�����j�E���   Q�l����j�U���   P�X����j�M���   R�D����j�E���   Q�0����j�U���   P�����j�M���   R�����j�E���   Q������j�U���   P������j�M���   R������j�E���   Q�����j�U���   P�����j�M���   R�����j�E���   Q�|����j�U���   P�h����j�M���   R�T����j�E���   Q�@����j�U���   P�,����j�M���   R�����j�E���   Q�����j�U���   P������j�M���   R������j�E���   Q������j�U���   P�����j�M���   R�����j�E���   Q�����j�U���   P�x����j�M���   R�d����j�E���   Q�P����j�U��   P�<����j�M��  R�(����j�E��  Q�����j�U��  P� ����j�M��  R������j�E��  Q������j�U��  P������j�M��  R�����j�E��   Q�����j�U��$  P�����j�M��(  R�t����j�E��,  Q�`����j�U��0  P�L����j�M��4  R�8����j�E��8  Q�$����j�U��<  P�����j�M��@  R������j�E��D  Q������j�U��H  P������j�M��L  R������j�E��P  Q�����j�U��T  P�����j�M��X  R�����j�E��\  Q�p����j�U��`  P�\����]�������̋�U��} u�   �E�;ȼtj�U�P�&�����M�Q;̼tj�E�HQ������U�B;мtj�M�QR�������E�H0;��tj�U�B0P�������M�Q4;��tj�E�H4Q�����]�����̋�U��} u�  �E�H;Լtj�U�BP�t�����M�Q;ؼtj�E�HQ�U�����U�B;ܼtj�M�QR�6�����E�H;�tj�U�BP������M�Q;�tj�E�HQ�������U�B ;�tj�M�Q R�������E�H$;�tj�U�B$P������M�Q8; �tj�E�H8Q������U�B<;�tj�M�Q<R�|�����E�H@;�tj�U�B@P�]�����M�QD;�tj�E�HDQ�>�����U�BH;�tj�M�QHR������E�HL;�tj�U�BLP� ����]�����������̋�U����EP�M������M(Q�U$R�E P�MQ�UR�EP�MQ�UR�M�����P�   ��$�E�M�����E��]���������̋�U��� �} ~,�EP�MQ�u  ���E�U�;U}�E���E��M�M�E�    �E�    �E�    �}$ u�U��H�M$j j �UR�EP3Ƀ}( ����   Q�U$R� �E��}� u3���  �}� ~63�u2�����3��u���r#h��  �M��T	R�.�����P�%������E���E�    �E�E�}� u3��  �M�Q�U�R�EP�MQj�U$R� ��u
�Y  �T  j j �E�P�M�Q�UR�EP�� �E��}� u
�,  �'  �M��   tI�}  t>�U�;U ~
�	  �  �E P�MQ�U�R�E�P�MQ�UR�� ��u
��   ��   ��   �E��E�}� ~63�u2�����3��u��r#h��  �U�DP�'�����P�������E���E�    �M��M��}� u�|�z�U�R�E�P�M�Q�U�R�EP�MQ�� ��u�V�T�}  u+j j j j �U�R�E�Pj �M$Q� �E��}� u�'�%�#j j �U R�EP�M�Q�U�Rj �E$P� �E��}� t�M�Q�������U�R�������E���]Ë�U����E�E��M�M��U��E����E���t�M����t�E����E��ۋE+E�����]����������̋�U����EP�M�����M$Q�U R�EP�MQ�UR�EP�MQ�M����P�"   �� �E�M��D���E��]�������������̋�U����E�    �} u�E��Q�Uj j �EP�MQ3҃}$ ��   R�EP� �E�}� u3��   3�u2�}� ~,�}����w#h��  �U�DP�4�����P�+������E���E�    �M�M��}� u3��a�U���Rj �E�P�{������M�Q�U�R�EP�MQj�UR� �E��}� t�EP�M�Q�U�R�EP�� �E��M�Q��������E���]�������̋�U���<�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� uh�?j jphx?j�=}������u̃}� u.詠���    j jphx?h�h�?�;���������R  �} t�} u	�E�    ��E�   �M̉MЃ}� uh0?j jshx?j��|������u̃}� u.�/����    j jshx?h�h0?������������   �}���v�E��@����	�M��U�Q�E��@B   �M��U�Q�E��M��UR�EP�MQ�U�R�U���E��} u�E��{�}� |X�E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj ��������Eă}��t�E���UU�B� �E��x }�����������]����������̋�U��� �E�����3��} ���E��}� u!hЇj h�   hx?j�g{������u̃}� u1�Ӟ���    j h�   hx?h��hЇ�b����������  �} t�} v	�E�   ��E�    �U�U�}� u!hp�j h�   hx?j��z������u̃}� u1�S����    j h�   hx?h��hp�����������d  �MQ�UR�EP�MQ�URhp���������E��}� }U�E�  �}�tI�}���t@�}v:�M��9��s����U��	�E���E�M�Qh�   �U��R�������}��uu3�t	�E�   ��E�    �M�M��}� u!h<�j h�   hx?j��y������u̃}� u.�V���� "   j h�   hx?h��h<�����������j�}� |a�}�t[�}���tR�E���;EsG�M����U+�9��s
����E���M����U+щU��E�Ph�   �M��U�D
P��������E���]���������������̋�U���,�E������E�    3��} ���E�}� u!hЇj h  hx?j��x������u̃}� u1�\����    j h  hx?h��hЇ����������  �} u�} u�} u3���  �} t�} v	�E�   ��E�    �U�U��}� u!hp�j h  hx?j�Wx������u̃}� u1�Û���    j h  hx?h��hp��R���������|  �M;M��   膛����U��EP�MQ�UR�E��P�MQhp��P������E��}��u~�}�t\�}���tS�U��;UsH�E���M+�9��s����U���E���M+ȉM�U�Rh�   �E�M�TR�����������8"u
�����M������  �`�Ϛ����U��EP�MQ�UR�EP�MQhp��������E��UU�B� �}��u"�}�u苚���8"u
聚���M������Y  �}� ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q�(������}��uu3�t	�E�   ��E�    �E܉E�}� u!h<�j hB  hx?j�Wv������u̃}� u.�Ù��� "   j hB  hx?h��h<��R�������������z�}�t\�}���tS�U���;UsH�E����M+�9��s����U���E����M+ȉM؋U�Rh�   �E��M�TR�F������}� }	�E�������E��EԋEԋ�]�������̋�U��EPj �MQ�UR�EP�MQ�@�����]�����������̋�U����EP�M������M������U���   �P�� �  �M�M�����E��]������������̋�U��j �EP������]�����������̋�U��j�h�h � d�    P��SVW�t�1E�3�P�E�d�    �=ص �tAj�{�����E�    h �hص�2������ص�E������   �j��{����ËM�d�    Y_^[��]����������������W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����������������̋�U�����}��E�P�   ���E��M#M�U��#U�ʉM�E�;E�t'�M�Q��  ��f�E��m���}��U�R�X   ���E�=�� tB�EP�MQ��  ���E�U�#���E�#��;�t�E�E�   ����E�E����E��]Ë�U����E�    �E��t	�M����M��U��t	�E����E��M��t	�U����U��E��t	�M����M��U�� t	�E����E��M��t�U���   �U��E%   �E��}�   �}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��   �U�t*�}�   t�}�   t�"�E��E���M���   �M���U���   �U��E%   t�M���   �M��E���]������̋�U���3�f�E��M��t�U���f�U��E��t�M���f�M��U��t�E���f�E��M��t�U���f�U��E��t�M��� f�M��U��   t�E���f�E��M��   �M��}�   w�}�   t&�}� t�}�   t&�B�}�   t+�7f�U�f�U��-�E�   f�E���M���   f�M���U���   f�U��E%   �E�t�}�   t�}�   t"�(�M���   f�M���U���   f�U��f�E�f�E��M��   t�U���   f�U�f�E���]��̋�U����E%�E�]��M�Q�`   ���E�U#U�E��#E�ЉU��M�;M�u�E��+�U�R�  ���E��E�P��\�����]��M�Q�   ����]�����������̋�U����E�    �E%�   t	�M����M��U��   t	�E����E��M��   t	�U����U��E%   t	�M����M��U��   t	�E����E��M��   t�U���   �U��E% `  �E��}� @  w�}� @  t$�}� t�}�    t#�:�}� `  t%�/�M��M��'�U���   �U���E�   �E���M���   �M��U��@�  �U�}�@t!�}� �  t&�}�@�  t�'�E�   �E���M���   �M���U���   �U��E���]������������̋�U����E�    �E��t�M��ɀ   �M��U��t�E�   �E��M��t�U���   �U��E��t�M���   �M��U��t�E�   �E��M��   t�U���   �U��E%   �E��}�   w�}�   t$�}� t�}�   t#�:�}�   t%�/�M��M��'�U��� @  �U���E�    �E���M��� `  �M��U��   �U�}�   t�}�   t�}�   t�$�E�@�  �E���M���@�M���U��� �  �U��E���]������������̋�U��h(��EP�MQ�	   ��]����̋�U���<�t�3ŉE�E�H
���  ���?  �M�U�B
% �  �E�M�Q�U܋E�H�M��U����E�}����u8�E�    �M�Q��  ����t	�E�    ��U�R�  ���E�   �Z  �E�P�M�Q�  ���U�U؋E�HQ�U�R�  ����t	�E���E�M�U�A+B9E�}�M�Q�*  ���E�    �E�   ��   �U�E�;Bk�M�Q�U�R�  ���E؉E�M�Q+U�UċE�P�M�Q�Z  ���U�BP�M�Q�  ���U�B��P�M�Q�1  ���E�    �E�   �~�U�E�;|B�M�Q�  ���U܁�   ��U܋E�HQ�U�R��  ���E��UJ�M��E�   �2�E�M�H�M��U܁�����U܋E�HQ�U�R�  ���E�    �E�H���    +щU��E��M���E܋M���Ɂ�   ���EԋU�z@u�E�MԉH�U�E����M�y u�U�Eԉ�E��M�3��������]��̋�U����E�    �E���E��M����M�E虃�����E�U��  �yJ���B�   +E�   �M���U��E�M��#U�t'�E�P�MQ�n   ����u�U�R�EP��   ���E�����M���E�M#��E�M���U���U��	�E���E�}�}�M�U��    ��E���]����������̋�U����E�������E��E%  �yH���@�   +ȉM����M����҉U��E��M��#U�t3��1�E����E��	�M����M��}�}�U��E�<� t3���߸   ��]������������̋�U����E�������E��E%  �yH���@�   +ȉM�   �M���U�E��M��R�E�P�M��U��P�V   ���E��M����M��	�U����U��}� |)�}� t#�E��M��Rj�E��M��R�   ���E��ȋE���]������̋�U����E�    �EE�E��M�;Mr�U�;Us	�E����E��M�U���E���]Ë�U����E�E��M�M��E�    �	�U����U��}�}�E�M����E���E�M����M��Ӌ�]��̋�U��Q�E�    �	�E����E��}�}�M��U��    ���]���������������̋�U��Q�E�    �	�E����E��}�}�M��U�<� t3���߸   ��]�������̋�U���V�E�������E��E%  �yH���@�E����M����҉U��E�    �E�    �	�E����E��}�}M�M��U��#E�E�M��U���M���M��U���E��M��U��E��M���    +M�U���U���E�   �	�E����E��}� |.�M�;M�|�U�+U��E��M�u������E��M��    ��^��]��̋�U��h@��EP�MQ�i�����]����̋�U���   �t�3ŉEčE��E�3�f�M��E�   �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    �E�    3҃}$ �U��}� u!h@�j h�   h��j�he������u̃}� u0�Ԉ���    j h�   h��h��h@��cq����3��  �M�M��U��U��	�E����E��M���� t!�E����	t�U����
t�M����u�Ƀ}�
�s  �E���M��U����U��E���x�����x����G  ��x����$��r�U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �`�M���t�����t���+t��t���-t#��t���0t�*�E�   �1�E�   3�f�U��"�E�   � �  f�E���E�
   �M����M��  �E�   �U���1|�E���9�E�   �M����M��   �U��E$����   ��;�u	�E�   �j�M���p�����p�����+��p�����p���:w8��p�����s�$�s�E�   �+�E�   �"�U����U��E�   ��E�
   �E����E���  �M���1|�U���9�E�   �E����E��K�M��U$����   ��;�u	�E�   �*�E���l�����l���0t�	�E�   ��E�
   �M��M��[  �E�   ��U���E��M����M��U���0|:�E���91�}�s �Mԃ��M��U���0�E���M����M��	�U����U���E��M$����   ��
;�u	�E�   �a�U���h�����h�����+��h�����h���:w/��h�����\s�$�Ps�E�   �"�E����E��E�   ��E�
   �M����M��w  �E�   �E�   �}� u'��U���E��M����M��U���0u�E����E�����M���U��E����E��M���0|8�U���9/�}�s'�Eԃ��E��M���0�U��
�E����E��M����M���U���d�����d�����+��d�����d���:w/��d������s�$��s�E�   �"�E����E��E�   ��E�
   �M����M��  �E�   �U���0|�E���9�E�   �M����M���E�
   �U��U��E  �E����E��M���1|�U���9�E�	   �E����E��U�M���`�����`���+t-��`���-t��`���0t�"�E�   �&�E�   �E�������E�   ��E�
   �U��U��  �E�   ��E���M��U����U��E���0u���M���1|�U���9�E�	   �E����E���E�
   �M����M��`  �U���1|�E���9�E�	   �M����M��*�U���\�����\���0t�	�E�   ��E�
   �E��E��  �E�   ǅ|���    ��M���U��E����E��M���0|:�U���91��|���k�
�M��TЉ�|�����|���P  ~ǅ|���Q  �묋�|����E���M���U��E����E��M���0|�U���9���E�
   �E����E��d�}  tN�M����M��U���X�����X���+t��X���-t��E�   �E�������E�   ��E�
   �E��E���E�
   �M����M������U�E���}� �9  �}� �/  �}� �%  �}�v+�M���|	�U����U��E�   �E����E��M����M��}� ��   �U����U��	�E����E��M����u�Eԃ��EԋM����M��ٍU�R�E�P�M�Q�#t  ���}� }�U��ډU��E�E��E��}� u	�M�M�M��}� u	�U�+U�U��}�P  ~	�E�   �B�}�����}	�E�   �0�EP�M�Q�U�R�  ��f�E�f�E�M��M�U��U�f�E�f�E��3�f�M�3�f�U��E�E؋M؉M�}� u$3�f�U�3�f�E��M�M؋U؉U�E܃��E��V�}� t(��  f�M��E�   ��E�    3�f�U�E܃��E��(�}� t"3�f�M�3�f�U��E�E؋M؉M�U܃��U܋Ef�M�f��U�E�B�M�U؉Q�E��M���Uf�B
�E܋M�3�������]Ë��j7k�kilMmBnndoo�o�p`p�k�k�k�k  �&mm8m  �nn-n  ̋�U����t�3ŉE��0���`�E��} u�   �} }�M�ىM�����`�U��} u3��Mf��} tr�U���T�U��E���E�M���M�}� u�׋U�k�U��U�E���� �  |#�U��E�J�M��R�U�E���E�M�M�U�R�EP�   ��눋M�3�������]�����������̋�U���L�t�3ŉE�3�f�E��E�    �E�    �E�    �E�    �Mf�Q
f�U�Ef�H
f�M��U��E�3Ё� �  f�U��M���  f�M��UЁ��  f�U��E��M��f�E��U���  }�E�=�  }�M�����  ~2�U���ҁ�   ��� ���E�P�M�A    �U�    �  �E�=�?  "�M�A    �U�B    �E�     ��  �M��u9f�U�f��f�U��E�H�����u�U�z u�E�8 u3ɋUf�J
�  �EЅ�uLf�M�f��f�M��U�B%���u3�M�y u*�U�: u"�E�@    �M�A    �U�    �I  �E�    �E�    �	�E����E��}���   �M���M��E�   �   +U��U��	�Eȃ��Eȃ}� ~x�MM��MċUỦU��E�L؉M��U���M���E��E�P�M�Q�U��P�"������E��}� t�M�f�T�f���E�f�T܋M����M��Ũ��U��y����E���E��<����M����?  f�M��U���~$�E�%   �u�M�Q�d  ��f�U�f��f�U����E���Qf�M�f��f�M��U���},�E؃�t	�Mԃ��MԍU�R�  ��f�E�f��f�E��̃}� t�M؃�f�M��U؁� �  �E�%�� = � u_�}��uP�E�    �}��u8�E�    �M����  u� �  f�U�f�E�f��f�E��f�M�f��f�M��	�Uރ��U��	�Eڃ��E��M����  |/�U���ҁ�   ��� ���E�P�M�A    �U�    �-�Ef�M�f��U�E܉B�M�U��Q�E��M���Uf�B
�M�3�������]����������̋�U����E���   �����ىM��U�B%   �����؉E��M���E��M�Q��U��E�P�M�Q��U��E�P��]��������������̋�U����E�H����Ɂ�   ��M��U�B�����%   ��E��M�Q��E�P�M�Q��U��E�P�M���U��E���]�����������̋�U���x�t�3ŉE��M  f�E��M   f�M���   f�U��E��C�E���E���E���E���E���E���E���E���E���E���E���E�?�E�   f�Ef�E�M�M؋U�U��E�% �  f�E��M���  f�M��U���t	�E�@-��M�A �U��uM�}� uG�}� uA3��Mf��U��� �  ��҃���-�E�P�M�A�U�B0�E�@ �   �  �M���  �e  �   �Ef��}�   �u�}� tP�M؁�   @uEj j|h��h��hX�hL�j�U��R�[����P�E������E�@�E�    ��   �M���tW�}�   �uN�}� uHj h�   h��h��h�h��j�U��R�?[����P��������E�@�E�    �   �}�   �uK�}� uEj h�   h��h��h��h��j�M��Q��Z����P�������U�B�E�    �Cj h�   h��h��hh�h`�j�E��P�Z����P�J������M�A�E�    �  �U���f�U��E�%�   f�E��M���f�M��U��E����M��E�����M��E����+U��U��M���f�M�f�U�f�U��E؉E��M��M�3�f�U�j�E���P�M�Q�A������U����?  |f�E�f��f�E��M�Q�U�R��������Ef�M�f��U��tP�E�E�E�} @3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �  �}~�E   �U����?  �U�3�f�E��E�    �	�M���M�}�}�U�R�S�������}� },�E���%�   �E��	�M����M��}� ~�U�R��������E���E��M���M��	�U���U�}� ~a�E��E̋M��MЋU��UԍE�P��������M�Q��������U�R�E�P�R  ���M�Q�������U���0�E���M����M��E� 됋U����U��E���M�U����U��E��5|[�	�M����M��U��9U�r�E����9u�U��0�ًE��9E�s�M����M��Uf�f���Mf��U���M���k�	�U����U��E��9E�r�M����0u�ߋE��9E�s=3ɋUf�
�E�- �  �������-�M�A�U�B�E�@0�M�A �   �&�U���E�+��M�A�U�B�M�D �E܋M�3�菸����]�����������̋�U����EP�M�R�E�Q�������E��}� t0�U��Rj�E�HQ�������E��}� t�U�B���M�A�U��R�E�HQ�U�BP�M������E�}� t�M�Q���E�P�M��Q�U�BP�M�QR��������]�̋�U��j�h8�h � d�    P���SVW�t�1E�3�P�E�d�    �E������E������}�u!�r���     �Zr��� 	   ��������  �} |�E;��s	�E�   ��E�    �MԉM܃}� uhp�j jMh�j�N������u̃}� u<�#r���     ��q��� 	   j jMh�h��hp��zZ�����������C  �E���M���������D
������؉E�uhċj jNh�j��M������u̃}� u<�q���     �_q��� 	   j jNh�h��hċ��Y�����������   �UR��g  ���E�    �E���M���������D
��t �MQ�UR�EP�MQ�   ���E��U��F��p��� 	   � q���     �E������E�����3�uh0�j jYh�j�#M������u��E������   ��MQ�#h  ��ËE��U�M�d�    Y_^[��]�������̋�U����E�E��M�M��UR�se  ���E�}��u;�2p��� 	   3�u!h0�j h�   h�j�L������u̃������   �UR�E�P�M�Q�U�R� !�E��}��u#�D �E��}� t�E�P�o�����������>�M���U���������L����U���E���������L�E��U���]��������̋�U��j�hX�h � d�    P���SVW�t�1E�3�P�E�d�    �}�u�co���     �(o��� 	   ����  �} |�E;��s	�E�   ��E�    �M؉M��}� uhp�j jCh��j�XK������u̃}� u9��n���     �n��� 	   j jCh��hЌhp��KW��������/  �E���M���������D
������؉E�uhċj jDh��j��J������u̃}� u9�nn���     �3n��� 	   j jDh��hЌhċ��V��������   �UR�d  ���E�    �E���M���������D
��t�MQ�UR�EP�   ���E��?�m��� 	   ��m���     �E�����3�uh0�j jOh��j�J������u��E������   ��EP�e  ��ËE�M�d�    Y_^[��]���������������̋�U�츐<  職���t�3ŉE��E�    �E�    �E�    �E��E�} u3���
  3Ƀ} ���M��}� uh��j jmh��j�XI������u̃}� u9��l���     �l���    j jmh��h��h���KU��������
  �E���M���������D
$�����E��M���t	�U���uo�E��������E�uhx�j juh��j�H������u̃}� u9�Rl���     �l���    j juh��h��hx��T���������	  �U���E���������T�� tjj j �EP�_������MQ�
  ����td�U���E���������T��   tA�����EԋEԋHl3҃y �U�E�P�M���U���������Q�!�E�}� ��  �}� t�U�����  �!�E��E�    �E�    �E�EЋM�+M;M�}  �U�����  �E��3҃�
�U��E���M���������|
8 ��   �E���M���������D
4P��������u!h@�j h�   h��j�G������u̋U���E���������T4�U��EЊ�M��U���E���������D8    j�U�R�E�P�gd  �����u�  �   �M��R�y���������   �E�+E�M+ȃ�v'j�U�R�E�P�d  �����u�O  �MЃ��M��K�U���E���������UЊ�T4�E���M���������D
8   �E����E���  �j�M�Q�U�R�c  �����u��  �EЃ��E��4�M���t	�U���u"�E�f�f�M��U�3���
���E��MЃ��M��U�����   j j j�E�Pj�M�Qj �U�R� �Eȃ}� u�f  �[j �E�P�M�Q�U�R�E���M���������
P�� ��t�M�+MM�M��U�;U�}�  ��D �E��	  �}� tl�E�   �E�j �E�P�M�Q�U�R�E���M���������
P�� ��t!�M�;M�}�   �U���U�E����E���D �E��   �   �M���t	�U���u{�E�P��_  �����U�;�u�E����E���D �E��R�}� tG�E�   �   f�M��U�R�_  �����M�;�u�U����U��E���E���D �E���t�����  �M���U���������L��   �k  �E�    �U����?  ǅ����    ǅ����    �E������������+M;M�  ������������������������+�=�  sz������+U;Usl�����������������������������������
u!�M���M싕�����������������������������������������������q���j �M�Q������������+�R������Q�U���E���������R�� ��t �E�E��E�������������+�9M�}���D �E��������  �E����C  �M������ǅ����    ������+U;U�  ������������������������+ʁ��  ��   ������+E;Esu������f�f����������������������������
u&�U���U�   ������f���������������������f������f����������������c���j �E�P������������+�Q������P�M���U���������Q�� ��t �U�U��U�������������+�9E�}���D �E���������  �U������ǅ����    �E������������+M;M��  ǅt���    ������������������������+�=�  sz������+U;Usl������f�f����������������������������
u�   ������f�
��������������������f������f����������������q���j j hU  ��x���Q������������++���P������Pj h��  � ��t�����t��� u�D �E��   �   ǅp���    j �M�Q��t���+�p���R��p�����x���Q�U���E���������R�� ��t��p���E���p�����D �E����t���;�p������t���;�p���~�������+E�E��U����Jj �M�Q�UR�EP�M���U���������Q�� ��t�E�    �U��U��	�D �E�}� ��   �}� t0�}�u�b��� 	   �b���M���U�R�a��������V�L�E���M���������D
��@t�M���u3��%��,b���    �Qb���     ������E�+E�M�3��$�����]Ë�U����} uh�kj j.h�j�]>������u̋T����T��U�U�j:hԍjh   茻�����E��E��M��H�}� t�U��B���M��A�U��B   �%�E��H���U��J�E����M��A�U��B   �E��M��Q��E��@    ��]��������������̋�U����}�u�a��� 	   3��   �} |�E;��s	�E�   ��E�    �M��M��}� uhp�j j(h��j�N=������u̃}� u*�`��� 	   j j(h��hl�hp��LI����3���E���M���������D
��@��]���̋�U��X�]����̋�U��Q�=�� u���   ��=��}
���   h�   h��jj���P�I������d��=d� u?���   h�   h��jj���Q�������d��=d� u
�   �   �E�    �	�U����U��}�}�E���X��M��d������E�    �	�E����E��}�}f�M����U����������<�t8�M����U����������<�t�M����U����������< u�M���ǁh������3���]����̋�U���[  �����t�VY  j�d�Q������]���̋�U��}X�r4�}��w+�E-X�����P�EB�����M�Q�� �  �E�P��M�� Q�� ]���������������̋�U��}}#�E��P��A�����M�Q�� �  �E�P��M�� Q�� ]���̋�U��}X�r4�}��w+�E�H������U�J�E-X�����P��A������M�� Q�� ]���������������̋�U��}}#�E�H������U�J�E��P�A������M�� Q�� ]���̋�U��Q3��} ���E��}� uh(nj j)h �j��9������u̃}� u+�_]���    j j)h �h�h(n��E���������U�B��]���������������̋�U��t���3�9X�����]����̋�U���@�} u�} v�} t	�E�     3���  �} t	�M���������;U����E�uh��j jJh��j� 9������u̃}� u0�\���    j jJh��h��h���E�����   �\  �UR�M������M������ �x ��   �M���   ~C�} t�} v�URj �EP�*������\��� *   �\����M؍M��
����E���  �} tw3�;U��؉E�uhx<j j]h��j�I8������u̃}� u=�[��� "   j j]h��h��hx<�GD�����E�"   �M������E��x  �U�E��} t	�M�   �E�    �M��g����E��J  �=  �E�    �U�Rj �EP�MQj�URj �M��e���� �HQ� �E��}� t
�}� ��   �}� ��   �D ��z��   �} t�} v�URj �EP������3�t	�E�   ��E�    �U��U܃}� uh<�j j{h��j�7������u̃}� u:�Z��� "   j j{h��h��h<��C�����E�"   �M��f����E��L�LZ��� *   �AZ����MȍM��D����E��*�} t�U�E���E�    �M��"����E���M�������]�̋�U��j �EP�MQ�UR�EP�������]��������������̋�U���L�E�    �} t�} u3��(  �} t�} v3��Mf�3҃} �U�}� uh��j jEhP�j��5������u̃}� u.�_Y���    j jEhP�h(�h����A��������  �MQ�M��Z����} �  �M��X�����z uj�E�;EsG�MM�f��Ef��MM����u�E��E؍M�������E��O  �M����M��U���U뱋E��EԍM�������E��%  �  �MQ�URj��EPj	�M��������QR� �E��}� t�E����EЍM��x����E���  �D ��zt*�PX��� *   3ɋUf�
�E������M��C����E��  �E�E��M�M��	�U���U�E��M����M���tk�U����ta�M��2���P�M��R��������t@�E��H��u,��W��� *   3ҋEf��E������M�������E��#  �	�M���M��|����U�+U�U܋EP�MQ�U�R�EPj�M�������QR� �E��}� u*�\W��� *   3��Mf��E������M��O����E��   �U��U��M��9����E��   �   �M��T���� �x u�MQ��=�����E��M������E��j�`j j j��URj	�M������ �HQ� �E��}� u!��V��� *   �E������M������E�� ��U����U��M������E���M�������]��̋�U���L�E�    �} u�} t�} t�} w	�E�    ��E�   �EĉE��}� u!h@�j h�   hP�j�2������u̃}� u3�V���    j h�   hP�h$�h@��>�����   ��  �} tY3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���E��M���Qh�   �U��R藜�����} t	�E�     �MQ�M������U;Uv�E�E���M�M��U��U�����;E�Ƀ��M�u!h��j h  hP�j�1������u̃}� u@�U���    j h  hP�h$�h���=�����E�   �M�������E���  �M�����P�E�P�MQ�UR��������E�}��ux�} tX3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P�c������KT����MЍM��N����E��/  �U���U�} ��   �E�;E��   �}���   3ɋUf�
�}�tK�}���tB�}v<�E��9��s����M��	�U���U��E���Ph�   �M��Q�ǚ�����U�9U����E�u!hȐj h  hP�j�0������u̃}� u=�xS��� "   j h  hP�h$�hȐ�<�����E�"   �M��U����E��9�U�U��E�P   3��M�Uf�DJ��} t�E�M��U��UȍM������Eȋ�]���̋�U��j �EP�MQ�UR�EP�MQ�`�����]�����������̋�U���4�} t�} v	�E�   ��E�    �E�E�}� uhYj jh(pj�/������u̃}� u0�wR���    j jh(phБhY�	;�����   �K  �} ��   �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q� �����3҃} �U��}� uhdXj jh(pj�F.������u̃}� u0�Q���    j jh(phБhdX�D:�����   �  �M�M��U�U��}� v�E����t�U����U��E����E��܃}� ��   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���M܋U�Rh�   �E��P��������o��t3�t	�E�   ��E�    �E؉E�}� uh�oj j h(pj�;-������u̃}� u0�P���    j j h(phБh�o�99�����   �{  �U��E��
�U���M����M��U���U��t�E����E�t�̓}� ��   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���MԋU�Rh�   �E��P��������<X��t3�t	�E�   ��E�    �EЉE�}� uh Xj j*h(pj�-,������u̃}� u-�O��� "   j j*h(phБh X�+8�����"   �p�}�th�}���t_�U+U���;UsQ�E+E����M+�9��s����U���E+E����M+ȉM̋U�Rh�   �E+E��M�TR������3���]�������������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�0   �E��j �MQ�UR�EP�MQ�   �E��E���]����������̋�U���03��} ���E�}� uh =j jfhВj��*������u̃}� u0�MN���    j jfhВh��h =��6�����   ��  3�;U��؉E�uh��j jghВj�*������u̃}� u0��M���    j jghВh��h���}6�����   �  �U� �}�tI�}���t@�}v:�E��9��s����M��	�U���UԋE�Ph�   �M��Q�~�����3҃} ��;U��؉E�uhH�j jihВj�)������u̃}� u0�*M��� "   j jihВh��hH��5�����"   ��  �}r�}$w	�E�   ��E�    �UЉU܃}� uh�j jjhВj�B)������u̃}� u0�L���    j jjhВh��h��@5�����   �O  �E�    �M�M��} t �U��-�E����E��M����M��U�ډU�E��E�E3��u�U�E3��u�E�}�	v�M��W�U��
�E����E���M��0�U��
�E����E��M����M��} v�U�;Ur��E�;Erl�M� �U�;U��؉E�u!h�j h�   hВj�8(������u̃}� u0�K��� "   j h�   hВh��h��34�����"   �E�U�� �E����E��M���U�E��M���E�M��U����U��E���E�M�;M�r�3���]� �������������̋�U���x�t�3ŉE��E�    �E�    �} t�} u3��  3��} ���EЃ}� uh��j jfhX�j�F'������u̃}� u.�J���    j jfhX�h,�h���D3��������8  �UR�M������} �.  �M������ �x ��   �M�;Msp�U�=�   ~"�EJ��� *   �E������M��@����E���  �MM��U���M��E���E��u�M��M��M��
����E��  �U����U�눋E��E��M�������E��  �  �M���������   ��   �} v�UR�EP�b  ���E�M�Qj �UR�EP�MQ�URj �M������ �HQ� �E��}� t3�}� u-�UU��B���u	�M����M��U��U��M��L����E���  �/I��� *   �E������M��*����E���  ��  �E�Pj �MQ�URj��EPj �M��/�����QR� �E��}� t�}� u�E����E��M��ӿ���E��j  �}� u�D ��zt"�H��� *   �E������M�蠿���E��7  �M�;M�  �U�Rj �M�访��� ���   Q�U�Rj�EPj �M�葿����QR� �E�}� t�}� t"�1H��� *   �E������M��,����E���  �}� |�}�v"�H��� *   �E������M�������E��  �E�E�;Ev�M��M��M��ݾ���E��t  �E�    ��U����U��E����E��M�;M�}4�UU��E��LԈ
�UU����u�M��M��M�舾���E��  벋U���U������E��E��M��b����E���   ��   �M��}�����y ur�E�    �U�U��	�Eȃ��EȋM����t;�E�����   ~"� G��� *   �E������M�������E��   �Ũ��U�벋ẺE��M��ڽ���E��t�j�M�Qj j j j��URj �M������ �HQ� �E��}� t�}� t�F��� *   �E������M�脽���E���U����U��M��n����E���M��a����M�3��g�����]���̋�U����E���E��M�M��U����U�t�E����t�U����U����}� t�E����u�E�+E������E��]�����̋�U���,�E�    �} t�} w�} u�} t	�E�    ��E�   �E�E��}� u!h �j h@  hX�j�"������u̃}� u3�qE���    j h@  hX�h�h �� .�����   �  �} tU�U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U��E�Ph�   �M��Q��������} t	�U�    �E;Ev�M�M���U�U܋E܉E�����;M�҃��U�u!h��j hL  hX�j�!������u̃}� u3�D���    j hL  hX�h�h���-�����   �  �MQ�U�R�EP�MQ�������E�}��ug�} tU�U� �}�tI�}���t@�}v:�E��9��s����M��	�U���U؋E�Ph�   �M��Q��������C��� �  �U���U�} ��   �E�;E��   �}���   �M� �}�tH�}���t?�}v9�U��9��s
����E��	�M���MԋU�Rh�   �E��P�_������M9M���ډU�u!hؓj hd  hX�j�������u̃}� u0�C��� "   j hd  hX�h�hؓ�+�����"   �(�M�M��E�P   �UU��B� �} t�E�M��E���]����������̋�U��j �EP�MQ�UR�EP�MQ������]�����������̋�U���D�E�    3��E܉E��E�E�E�E��E�M؉M�3҃} �Uԃ}� u!h�?j h�   hДj�������u̃}� u1�B���    j h�   hДh��h�?�*��������  �} t�} u	�E�    ��E�   �M̉MЃ}� u!h0?j h�   hДj�*������u̃}� u1�A���    j h�   hДh��h0?�%*��������8  �E��@B   �M��U�Q�E��M��}���?v�U��B�����E���M��A�UR�EP�MQ�U�R�U���E��} u�E���   �}� ��   �E��H���MȋU��EȉB�}� |!�M��� 3�%�   �EċM�����E����M�Qj �Wb�����Eă}��tY�U��B���E��M��U��Q�}� |"�E��� 3ҁ��   �U��E�����U��
��E�Pj �b�����E��}��t�E�� 3ɋU�Ef�LP��M��y }�����������]��������������̋�U���,�E������E�    3��} ���E�}� u!hЇj h9  hДj�`������u̃}� u1��?���    j h9  hДh|�hЇ�[(��������&  �} u�} u�} u3��  �} t�} v	�E�   ��E�    �U�U��}� u!h8�j h?  hДj��������u̃}� u1�3?���    j h?  hДh|�h8���'��������  �M;M��   ��>����U��EP�MQ�UR�E��P�MQh0��P������E��}����   �}�t^�}���tU�U��;UsJ�E���M+�9��s����U���E���M+ȉM�U���Rh�   �E�M�TAR�o������W>���8"u
�M>���M�������  �c�9>����U��EP�MQ�UR�EP�MQh0��������E�3ҋE�Mf�TA��}��u"�}�u��=���8"u
��=���U������a  �}� ��   3��Mf��}�tJ�}���tA�}v;�U��9��s
����E��	�M���M��U���Rh�   �E��P茄�����}��ux3�t	�E�   ��E�    �U܉U�}� u!h<�j hf  hДj�������u̃}� u1�'=��� "   j hf  hДh|�h<��%��������   ����|�}�t^�}���tU�M���;MsJ�U����E+�9��s����M���U����E+E؋M���Qh�   �U��E�LPQ襃�����}� }	�E�������U��UԋEԋ�]������̋�U��EPj �MQ�UR�EP�MQ�0�����]�����������̋�U��Q�E�    �}
u"�} }j�EP�MQ�UR�EP�0   �E��j �MQ�UR�EP�MQ�   �E��E���]����������̋�U���03��} ���E�}� uh =j jfhВj�1������u̃}� u0�;���    j jfhВh��h =�/$�����   �  3�;U��؉E�uh��j jghВj��������u̃}� u0�;;���    j jghВh��h����#�����   �  3ҋEf��}�tK�}���tB�}v<�M��9��s����U��	�E���EԋM���Qh�   �U��R�ʁ����3��} ����;E��ىM�uhH�j jihВj�
������u̃}� u0�v:��� "   j jihВh��hH��#�����"   ��  �}r�}$w	�E�   ��E�    �EЉE܃}� uh�j jjhВj�������u̃}� u0��9���    j jjhВh��h��"�����   �`  �E�    �U�U��} t%�-   �M�f��U����U��E����E��M�ىM�U��U�E3��u�U�E3��u�E�}�	v�E��W�M�f��U����U���E��0�M�f��U����U��E����E��} v�M�;Mr��U�;Urn3��Mf��U�;U��؉E�u!h�j h�   hВj�{������u̃}� u0��8��� "   j h�   hВh��h��v!�����"   �M3ҋE�f��M����M��U�f�f�E��M��U�f�f��M�f�U�f��E����E��M���M�U�;U�r�3���]� ��������̋�U����s�����   u<�E�8csm�t1�M�9&  �t&�U�%���="�r�M�Q ��t
�   ��   �E�H��ft4�U�z t�} uj��EP�MQ�UR��  ���   ��   �   �E�x u$�M��������!���   �E�x ��   �M�9csm�uX�U�zrO�E�x"�vC�M�Q�B�E��}� t1�M$Q�U R�EP�MQ�UR�EP�MQ�UR�U��� �E��E��0�)�E P�MQ�U$R�EP�MQ�UR�EP�MQ�   �� �   ��]�������������̋�U���D�E� �E� �E�x�   �M�Q���   �E��	�M�Q�U��E��E��}��|�M�U�;Q}���B���E�8csm��[  �M�y�N  �U�z �t�E�x!�t�M�y"��&  �U�z �  �s������    u��  �`������   �E�R������   �M�E�j�UR��J  ����t��<B���E�8csm�u;�M�yu2�U�z �t�E�x!�t�M�y"�u�U�z u��A���������    ty�ӌ�����   �E��Ō��ǀ�       �M�Q�UR�^  ������t�C�M�Q�  ���Ѕ�t+j�EP�4  ��h���M���  ht��M�Q�FJ  ��@���U�:csm��n  �E�x�a  �M�y �t�U�z!�t�E�x"��9  �M�y �+  �U�R�E�P�M�Q�U R�EP�Ń�����E���M����M��U���U�E�;E���   �M�;U��E�M�;H~�ˋU�B�E��M�Q�U���E���E�M����M��}� ��   �U�B�H���M؋U�B�H��U���E܃��E܋M؃��M؃}� ~d�U؋�EԋM�QR�E�P�M�Q��  ����u���E��U�R�E$P�M Q�U�R�E�P�M�Q�UR�EP�MQ�UR�EP�f  ��,�	���D���������M��tj�UR�  ���E�����   �M��������!���   �E�x ��   �M�QR�EP�=  ���ȅ���   �z������   �U��l������   �E��^����M���   �P����U���   �}$ u�EP�MQ�����UR�E$P��~��j��MQ�UR�EP�  ���M�QR�s  ��������M���   �����U���   �@�E�x v7�M��u*�U$R�E P�M�Q�UR�EP�MQ�UR�EP��   �� ��>��蝉�����    u��>����]���������̋�U��Q�M��EP�M���G  �M��ĕ�E���]� ��������̋�U��Q�M��E�� ĕ�M��vH  ��]��̋�U��Q�M��M�������E��t�M�Q��e�����E���]� �̋�U��Q�M��EP�M��G  �M��ĕ�E���]� ��������̋�U���V�E�8  �u�c  貈�����    tW褈�����݃��9��   tC�M�9MOC�t8�U�:RCC�t-�E$P�M Q�UR�EP�MQ�UR�EP�~������t��   �M�y t��R=���U�R�E�P�MQ�U R�EP�������E���M����M��U����U��E�;E���   �M��U;|\�E��M;HQ�U��B�����M��Q�| t�E��H�����U��B�L�Q��u�E��H�����U��B���@t�w���j�U$R�E P�M�Qj �U��B�����M�AP�UR�EP�MQ�UR�EP��  ��,�3���^��]���������������̋�U��Q�E�x t�M�Q�B��u
�   �   �M�U�A;Bt$�M�Q��R�E�H��Q袁������t3��O�U���t
�M���t1�E���t
�U���t�M���t
�E���t	�E�   ��E�    �E���]����̋�U����E��M��U���E��}�RCC�t(�}�MOC�t�}�csm�t�@�V���ǀ�       �:���B������    ~�4����   �E�M����E�3��3���]�����̋�U��j�hȢh � d�    P���SVW�t�1E�3�P�E�d�    �e�E�x�   �M�Q���   �E��	�M�Q�U܋E܉E�觅���   �E؋M؋���E؉�E�    �M�;M��   �}��~�U�E�;B}��w:���M�Q�E�M��E�   �U�B�M�|� t%�U�E��Bh  �MQ�U�B�M�T�R�l
  �E�    ��E�P�z�����Ëe��E�    �M��M��f����E������   �)�ބ�����    ~�Є���   �EԋUԋ���MԉËU�;Uu��9���E�M�H�M�d�    Y_^[��]Ë�U����E�E��}  t�M Q�UR�E�P�MQ�  ���}, u�UR�EP�!y����MQ�U,R�y���E$�Q�UR�EP�M�Q�������U$�B���M�Ah   �U(R�E�HQ�UR�EP�M�Q�UR�$   ���E��}� t�EP�M�Q�[x����]�������̋�U��j�h�h � d�    P���SVW�t�1E�3�P�E�d�    �e�E�E��E�    �M�Q��U��E�HQ�U�R��{�����E��j������   �E��\������   �M��N����U���   �@����M���   �E�    �E�   �E�   �U R�EP�MQ�UR�EP�yx�����E��E�    ��   �M�Q�  ��Ëe�����ǀ      �U�B�E��M�y�   �U�B%�   �ȉM��	�U�B�E��M��M��U�B�E��E�    �	�Mă��MċU�E�;BsG�M�k��U��E�;D
~3�M�k��U��E�;D
!�M�k��U��D
���E��M��U��ʉE��륋M�Q�URj �EP�������E�    �E�    �E������E�    �   �   �M�U��Q��E�P�z�����ށ���Mȉ��   �Ё���Ủ��   �E�8csm�u\�M�yuS�U�z �t�E�x!�t�M�y"�u/�}� u)�}� t#�U�BP��y������t�M�Q�UR�  ��ËEЋM�d�    Y_^[��]����������̋�U��Q�E��M��U��:csm�uN�E��xuE�M��y �t�U��z!�t�E��x"�u!�M��y u����ǀ     �   ��3���]���̋�U��j�h�h � d�    P���SVW�t�1E�3�P�E�d�    �e��E�    �E�x t#�M�Q�B��t�M�y u�U�%   �u3���  �M���   �t�E�E���M�Q�E�L�M��E�    �U���tXj�M�QR��=  ����t9j�E�P�=  ����t'�M��U�B��M��Q�U��P�G  ���M�����4���@  �U���txj�M�QR�k=  ����tYj�E�P�Y=  ����tG�M�QR�E�HQ�U�R�D�����E�xu"�M��9 t�U��R�E��Q��  ���U����f4���   �E�x uZj�M�QR��<  ����t>j�E�P��<  ����t,�M�QR�E��P�M�QR�g  ��P�E�P�
D������ 4���[j�M�QR�<  ����tAj�E�P�~<  ����t/�M�QR�k<  ����t�E���t	�E�   ��E�   ��3���E�������   Ëe���2���E������E�M�d�    Y_^[��]Ë�U��j�h8�h � d�    P���SVW�t�1E�3�P�E�d�    �e�E���   �t�U�U���E�H�U�D
�E��E�    �MQ�UR�EP�MQ�������E��}�t�}�t+�R�U��R�E�HQ�#  ��P�U�BP�M�Q�or���)j�U��R�E�HQ��   ��P�U�BP�M�Q�Dr���E�������   Ëe���1���E������M�d�    Y_^[��]����̋�U��j�hX�h � d�    P��SVW�t�1E�3�P�E�d�    �e�} t�E�8csm�t�U�M�y tL�U�B�x t@�E�    �M�Q�BP�M�QR�q���E�������E�����Ëe��1���E������M�d�    Y_^[��]�̋�U��Q�E�M�M��U�z |'�E�H�U�
�M�Q�M��M��U�E�B�E��E���]��������̋�U����} t��K1���} u�0���E� �E�    �	�E���E�M�U�;}m�E�H�Q���U��E�H�Q��E���M����M��U����U��}� ~4�E���M�U�BP�M�Q�U����EPR�t�������t�E���뀊E��]������������̋�U��j�h�d�    PQSVW�t�3�P�E�d�    �e��`{�����    u��`0���E�    �$0���$�={���M���   j j �9  �E����������E������r/���M�d�    Y_^[��]Ë�U��Q�E�    �	�E����E��M�U�;}'hؿ�E����M�Q�L��c������t����2���]��U���SQ�E���E��EU�u�M�m��t��VW��_^��]�MU���   u�   Q�t��]Y[�� ���̋�U���4  �t�3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M������E�    3Ƀ} �������������� u!h(nj h  h�mj�4�������u̃����� uF�"���    j h  h�mhԖh(n�,����ǅ��������M��w���������  �E�������������Q��@��   ������P�������������������t-�������t$����������������������������
ǅ�������������H$�����х�uV�������t-�������t$����������������������������
ǅ�������������B$�� ���ȅ�tǅ����    �
ǅ����   ������������������ u!h�lj h  h�mj��������u̃����� uF�(!���    j h  h�mhԖh�l�	����ǅ��������M�����������  3Ƀ} �������������� u!h�?j h  h�mj�7�������u̃����� uF� ���    j h  h�mhԖh�?�/	����ǅ��������M��z���������  ǅ����    �E�    ǅ����    �E�    �E�    �E��������������E���E���
  ������ ��  �������� |%��������x��������X����������
ǅ����    ������������������k�	��������x�����������������   3�tǅ����   �
ǅ����    ������������������ u!h0�j h`  h�mj���������u̃����� uF�4���    j h`  h�mhԖh0�������ǅ��������M�����������  ��������������������  �������$�|��E�    �M������P������R�Ѕ��������   ������P�MQ������R�]  ���E��������U���U����������؉�����u!h�lj h�  h�mj���������u̃����� uF�2���    j h�  h�mhԖh�l������ǅ��������M�����������  ������R�EP������Q�  ����  �E�    �UԉU؋E؉E�M�M��E�    �E������E�    �  �������������������� ������������wK�����������$����E����E��,�M����M��!�U����U���E��   �E��	�M����M��  ��������*u(�EP�tA�����E�}� }�M����M��U��ډU���E�k�
�������TЉU���  �E�    ��  ��������*u�MQ�A�����EЃ}� }�E�������U�k�
�������LЉM��  ��������������������I������������.�  �����������$����E���lu�U���U�E�   �E��	�M����M���   �U���6u&�M�Q��4u�E���E�M��� �  �M��   �U���3u#�M�Q��2u�E���E�M�������M��S�U���dt7�M���it,�E���ot!�U���ut�M���xt�E���Xu�ǅ����    ������U��� �U���E�   �E��D
  ��������������������A������������7�  ��������H��$���U���0  u�E�   �E��M���  tUǅ����    �UR�?����f������������Ph   ������Q�U�R������������������ t�E�   �&�EP��>����f��|�����|����������E�   �������U��W  �EP��>������x�����x��� t��x����y u����U��E�P������E��P�M���   t&��x����B�E���x�����+����E��E�   ��E�    ��x����B�E���x�����U���  �E�%0  u�M���   �M��}��uǅ��������	�UЉ�������������p����MQ��=�����E��U���  te�}� u����E��E�   �M���l�����p�����p�������p�����t��l������t��l�������l����ɋ�l���+M����M��[�}� u	����U��E���t�����p�����p�������p�����t��t������t��t�������t����ɋ�t���+E��E��  �MQ�=������h���肻������   3�tǅ����   �
ǅ����    ��������d�����d��� u!hXlj h�  h�mj���������u̃�d��� uF�<���    j h�  h�mhԖhXl�� ����ǅ��������M�����������  ��  �U��� t��h���f������f����h�����������E�   �  �E�   �������� �������U���@�U��������E��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Bh�  h$lj�UЁ�]  R�q�����E��}� t�E��E��MЁ�]  �M���EУ   �U���U�E�H��P���X�����\����M��'���P�E�P�M�Q������R�E�P�M�Q��X���R��P� �Ѓ��M���   t$�}� u�M��ݍ��P�U�R�$�P� �Ѓ���������gu*�U���   u�M�訍��P�E�P� �Q� �Ѓ��U����-u�M���   �M��U����U��E�P��������E��	  �M���@�M��E�
   �o�E�
   �f�E�   ǅ����   �
ǅ����'   �E�   �U���   t�E�0��������Q�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�	:������H�����L����   �U���   t�EP��9������H�����L����   �M��� tB�U���@t�EP�9��������H�����L�����MQ�x9���������H�����L����=�U���@t�EP�R9�������H�����L�����MQ�79����3҉�H�����L����E���@t@��L��� 7|	��H��� s,��H����ً�L����� �ډ�@�����D����E�   �E����H�����@�����L�����D����E�% �  u&�M���   u��@�����D����� ��@�����D����}� }	�E�   ��M�����M��}�   ~�E�   ��@����D���u�E�    �E��E��MЋUЃ��UЅ���@����D���t{�E��RP��D���Q��@���R��^����0��T����E��RP��D���P��@���Q�J^����@�����D�����T���9~��T����������T����E���T�����U����U��g����E�+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@t?�E�%   t�E�-�E�   �(�M���t�E�+�E�   ��U���t�E� �E�   �E�+E�+E䉅<����M���u������R�EP��<���Qj �  ��������R�EP�M�Q�U�R�8  ���E���t$�M���u������R�EP��<���Qj0��  ���}� ��   �}� ��   ǅ$���    �U���8����E܉�4�����4�����4�������4�������   ��8���f�f������������Rj��(���P��0���Q�Ϸ������$�����8�������8�����$��� u	��0��� uǅ���������&������P�MQ��0���R��(���P�;  ���Z����������Q�UR�E�P�M�Q�  �������� |$�U���t������P�MQ��<���Rj �  ���}� tj�E�P�Hw�����E�    ����������� t������tǅ����    �
ǅ����   �������� ����� ��� u!hЕj h�  h�mj�4�������u̃� ��� uC����    j h�  h�mhԖhЕ�,�����ǅ��������M��w����������������� ����M��[����� ����M�3��[U����]ÍI �����������#�^�a�l�V�K�y��� �I ��C�`�N�Y� ���������E��������������������   	
��U����E�H��@t�U�z u�E����U�
�s�E�H���M��U�E��B�}� |&�M��E��M���   �M��U����M���UR�EP�V0�����E��}��u�M�������U����M���]��������������̋�U��E�M���M��~!�UR�EP�MQ�)������U�:�u���]��������̋�U��Q�E�H��@t�U�z u�E�M�U�
�`�E�M���M��~P�U��E��MQ�UR�E�P�������M���M�U�:�u �����8*u�EP�MQj?��������렋�]����U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����t�3ŉE��N@  f�E��M�    �U�B    �E�@    ��M���M�U���U�} vt�E��M�P�U��@�E�MQ��������UR赒�����E�P�MQ�5������UR虒�����E��M��E�    �E�    �U�R�EP�������t����M�y uB�U�B���M�A�U�B���M���M�A�U����M��U���f�U�뵋E�H�� �  u�UR������f�E�f��f�E��؋Mf�U�f�Q
�M�3���P����]��������������̋�U��Q�} ��   �E;����   �M���U���������L����   �U���E���������<�th�=8�u<�U�U��}� t�}�t�}�t�"j j��!�j j��!�
j j��!�E���M�������������3�����
��� 	   ����     �����]������������̋�U����}�u��
���     �
��� 	   ����2  �} |�E;��s	�E�   ��E�    �M�M��}� u!hp�j h;  h�j���������u̃}� u<�{
���     �@
��� 	   j h;  h�h�hp������������   �E���M���������D
������؉E�u!hċj h<  h�j�S�������u̃}� u9��	���     �	��� 	   j h<  h�h�hċ�C����������U���E�����������]��������������̋�U��j�hУh � d�    P���SVW�t�1E�3�P�E�d�    �E���M��������M��E�   �U��z u_j
�������E�    �E��x u,h�  �M���Q�` ��u�E�    �U��B���M��A�E������   �j
�z�����Ã}� t!�U���E���������TR�� �E�M�d�    Y_^[��]����������̋�U��E���M���������D
P�� ]��������̋�U��Q�=���u�|  �=���u���  �(j �E�Pj�MQ���R�� ��u���  �f�E��]Ë�U���$�} t�} u3���  �E���u�} t3ҋEf�3���  �MQ�M���}���M���~������   t1�M��~��� ���   thؗj jGhx�j���������u̍M��~����z u*�} t�Ef��Uf�
�E�   �M��4~���E��R  �M��T~��P�E�Q�'n��������   �M��4~������   ~R�M��!~��� �M;��   |=3҃} ��R�EP�M���}������   R�EPj	�M���}����QR� ��uB�M���}��� �M;��   r�U�B��u"�r��� *   �E������M��m}���E��   �M��}������   �U�M��J}���E��k�a3��} ��P�MQj�URj	�M��U}��� �HQ� ��u� ��� *   �E������M���|���E���E�   �M���|���E���M���|����]������̋�U��j �EP�MQ�UR�������]���̋�U��j�h�h � d�    P���SVW�t�1E�3�P�E�d�    �E�    j��������E�    �E�   �	�E����E��M�;����   �U�d��<� t|�M��d����H��   t"�U�d���Q�  �����t	�U���U�}�|=�E��d����� R�l j�E��d���R��j�����E��d���    �Y����E������   �j�a�����ËE�M�d�    Y_^[��]��������̋�U��} uj �.  ���@�EP�@   ����t����+�M�Q�� @  t�EP荦����P��  ������3�]�������̋�U����E�    �E�E�M�Q����u|�E�H��  tn�U�E�
+H�M��}� ~Z�U�R�E�HQ�U�R������P�>�����;E�u�E�H��   t�U�B����M�A��U�B�� �M�A�E������U�E�H�
�U��B    �E���]�����̋�U��j�   ��]���������������̋�U��j�h�h � d�    P���SVW�t�1E�3�P�E�d�    �E�    �E�    j�y������E�    �E�    �	�E����E��M�;����   �U�d��<� ��   �M��d����H��   ��   �U�d���Q�U�R��������E�   �E��d����B%�   te�}u%�M��d���P����������t	�M���M��:�} u4�U�d����Q��t!�E��d���R���������u�E������E�    �   ��E��d���R�E�P�������������E������   �j������Ã}u�E����E܋M�d�    Y_^[��]���������������̋�U����  �t�3ŉE�ǅ����    �E�    �E�    �E�    �E�    �E�    �E�    �EP�M��[w���E�    3Ƀ} �������������� u!h(nj h  h�mj�t�������u̃����� uF�� ���    j h  h�mh��h(n�l�����ǅ@��������M��w����@�����  3��} �������������� u!h�?j h  h�mj���������u̃����� uF�U ���    j h  h�mh��h�?�������ǅ<��������M��/w����<����r  ǅ����    �E�    ǅ����    �E�    �E�    �Uf�f�������������U���U���`  ������ �S  �������� |%��������x��������X�����(����
ǅ(���    ��(���������������k�	��������x�����������������   3�tǅ$���   �
ǅ$���    ��$��������������� u!h0�j h`  h�mj�~�������u̃����� uF������    j h`  h�mh��h0��v�����ǅ8��������M���u����8����  �������� ����� ����"  �� ����$��E�   ������Q�UR������P��  ����  �E�    �MԉM؋U؉U�E�E��E�    �E������E�    �  ������������������ ����������wL�������T�$�<�U����U��-�E����E��"�M����M���U��ʀ   �U��	�E����E��E  ��������*u(�UR��!�����E�}� }�E����E��M��ىM���U�k�
�������LЉM���  �E�    ��  ��������*u�EP�!�����EЃ}� }�E�������M�k�
�������DЉE��  ������������������I����������.�  �������|�$�h�U���lu�M���M�U���   �U��	�E����E���   �M���6u%�E�H��4u�U���U�E� �  �E��   �M���3u"�E�H��2u�U���U�E�%����E��S�M���dt7�E���it,�U���ot!�M���ut�E���xt�U���Xu�ǅ����    �w�����M��� �M���U���   �U��n
  ������������������A����������7�J  ���������$���M���0  u	�U��� �U��E�   �EP������f�������M��� tW���������   ������ƅ���� �M��r��P�M��{r��� ���   Q������R������P�?�������}�E�   �f������f�������������U��E�   �  �EP�C���������������� t�������y u����U��E�P�������E��P�M���   t&�������B�E���������+����E��E�   ��E�    �������B�E���������U���  �E�%0  u	�M��� �M��}��uǅ�������	�UЉ����������������MQ�s�����E��U��� ��   �}� u����E��M��������E�    �	�U܃��U܋E�;�����}L���������t?�M���p��P�������Q��`������t������������������������������d�}� u	����M��E�   �U�����������������������������t���������t���������������ɋ�����+U����U��  �EP�m������|����ߛ������   3�tǅ���   �
ǅ���    �������x�����x��� u!hXlj h�  h�mj�0�������u̃�x��� uF�����    j h�  h�mh��hXl�(�����ǅ4��������M��so����4����  ��  �M��� t��|���f������f����|�����������E�   �  �E�   �������� f�������M���@�M��������U��E�   �}� }	�E�   �+�}� u��������gu	�E�   ��}�   ~�E�   �}У   ~Ah�  h$lj�MЁ�]  Q�pQ�����E��}� t�U��U��E�]  �E���EУ   �M���M�U�B��J���p�����t����M��n��P�U�R�E�P������Q�U�R�E�P��p���Q��R� �Ѓ��E�%�   t%�}� u�M��:n��P�M�Q�$�R� �Ѓ���������gu)�M���   u�M��n��P�U�R� �P� �Ѓ��M����-u�E�   �E��M����M��U�R�V������E��  �E���@�E��E�
   �u�E�
   �l�E�   ǅ����   �
ǅ����'   �E�   �M���   t�0   f�U싅������Qf�E��E�   ��E�   �M���   t�U���   �U��E�% �  t�MQ�a������`�����d����   �U���   t�EP�9������`�����d����   �M��� tB�U���@t�EP����������`�����d�����MQ�����������`�����d����=�U���@t�EP��������`�����d�����MQ�����3҉�`�����d����E���@t@��d��� 7|	��`��� s,��`����ً�d����� �ډ�X�����\����E�   �E����`�����X�����d�����\����E�% �  u&�M���   u��X�����\����� ��X�����\����}� }	�E�   ��M�����M��}�   ~�E�   ��X����\���u�E�    �������E��MЋUЃ��UЅ���X����\���t{�E��RP��\���Q��X���R�1?����0��l����E��RP��\���P��X���Q�>����X�����\�����l���9~��l����������l����E���l�����U����U��g���������+E��E܋M����M��U���   t)�}� t�E����0t�U����U��E�� 0�M܃��M܃}� ��  �U���@tN�E�%   t�-   f�M��E�   �2�U���t�+   f�E��E�   ��M���t�    f�U��E�   �E�+E�+E䉅T����M���u������R�EP��T���Qj �  ��������R�EP�M�Q�U�R��  ���E���t$�M���u������R�EP��T���Qj0�_  ���}� ��   �}� ��   �U���P����E܉�L�����L�����L�������L�����~}�M��i��P�M��|i��� ���   Q��P���R������P�@�������H�����H��� ǅ���������2������Q�UR������P�Z  ����P����H�����P����j����������R�EP�M�Q�U�R��  �������� |$�E���t������Q�UR��T���Pj �Y  ���}� tj�M�Q�W�����E�    �{��������� t������tǅ���    �
ǅ���   �������D�����D��� u!hЕj h�  h�mj��������u̃�D��� uC������    j h�  h�mh��hЕ������ǅ0��������M���g����0������������,����M��g����,����M�3��5����]�0�W��� �M�Y����������������� �I 	��������� ����Z�W�����(�5�����P�m�G�c�J�   	
��U��E�H��@t�U�z u�E����U�
�4�EP�MQ��   ���Ё���  u�E� ������M����E�]��̋�U��E�M���M��~!�UR�EP�MQ�y������U�:�u���]��������̋�U��Q�E�H��@t�U�z u�E�M�U�
�b�E�M���M��~R�Uf�f�E��MQ�UR�E�P�������M���M�U�:�u �����8*u�EP�MQj?���������랋�]�̋�U���8�t�3ŉE�V�E�H��@�d  �UR蕐�������t@�EP脐�������t/�MQ�s����������UR�b�������������E���E����E�H$�����у�tj�EP�+��������t@�MQ���������t/�UR�	����������EP���������������E���E����M�Q$������uh�M�Q���U��E�M��H�}� |2�U�f�Mf��U����  f�UދE����U�
f�E��  ��EP�MQ��  ���  �(  �UR�Y��������t@�EP�H��������t/�MQ�7����������UR�&�������������E���E����E��H��   ��   �URj�E�P�M�Q胒������t
���  ��   �E�    �	�U����U��E�;E�}s�M�Q���UԋE�MԉH�}� |.�U��M��T��E�����   �UЋE����U�
��EP�M��T�R������EЃ}��u���  �k�|����E%��  �[�E�H���M̋U�ẺB�}� |/�M�f�Ef��M����  f�MʋU����M�f�E����UR�EP�r  ��^�M�3��0����]ËD$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� �����������̋�U��Q�E�   �} u�E�    �E���]���������������̋�U��� VW�   ���}��E�E��M�M��} t�U���t�E� @��M�Q�U�R�E�P�M�Q� _^��]� �����̋�U��Q�M��M���   �E��t�M�Q������E���]� �̋�U��Q�M��E�� ��M��A    �U��B �E�Q�M���   �E���]� �����̋�U��Q�M��E�� ��M��A    �U��B �EP�M��   �E���]� �������̋�U��Q�M��E�;Et0�M���   �M�Q��t�E�HQ�M��m   ��U��E�H�J�E���]� �����̋�U��Q�M��E�� ��M��   ��]��̋�U����M��E��x t�M��Q�U���E���E���]���̋�U����M��} tK�EP���������E��M�Q�0�����U��B�E��x t�MQ�U�R�E��HQ��������U��B��]� �������������̋�U��Q�M��E��H��t�U��BP�0�����M��A    �U��B ��]��������̋�U��j j jj jh   @h$��!���]����������̋�U��=���t�=���t���P�!]�����������̋�U��j�h8�h � d�    P���SVW�t�1E�3�P�E�d�    �E�����3��} ���E��}� uh(nj j.hH�j�`�������u̃}� u+������    j j.hH�h4�h(n�^���������W�U�B��@t�M�A    �=�UR覈�����E�    �EP�C   ���E��E������   ��MQ������ËE�M�d�    Y_^[��]�������������̋�U����E�����3��} ���E�}� uhȘj jYhH�j�z�������u̃}� u.������    j jYhH�h��hȘ�x���������   �U�U��E��H��   ta�U�R�������E��E�P�  ���M�Q������P�  ����}	�E������$�U��z tj�E��HQ�L�����U��B    �E��@    �E���]�������̋�U��j�hX�h � d�    P���SVW�t�1E�3�P�E�d�    �}�u������ 	   ����  �} |�E;��s	�E�   ��E�    �M؉M��}� uhp�j j,h�j�#�������u̃}� u.����� 	   j j,h�h �hp��!���������;  �E���M���������D
������؉E�uhșj j-h�j��������u̃}� u.����� 	   j j-h�h �hș�����������   �UR�������E�    �E���M���������D
��t;�MQ�������P�!��u�D �E���E�    �}� u�>�����U��x���� 	   �E�����3�uh0�j jEh�j���������u��E������   ��UR�������ËE�M�d�    Y_^[��]���������̋�U��� �} uh�kj jdh0kj�m�������u̋M�M��U�R�5������E��E��H��   u&����� 	   �U��B�� �M��A���  �c  �/�U��B��@t$����� "   �M��Q�� �E��P���  �2  �M��Q��tJ�E��@    �M��Q��t�E��M��Q��E��H����U��J��E��H�� �U��J���  ��  �E��H���U��J�E��H���U��J�E��@    �E�    �M��M�U��B%  u6�`����� 9E�t�S�����@9E�u�M�Q肁������u�U�R袀�����E��H��  �  �U��E��
+Hy!h�jj h�   h0kj��������u̋E��M��+Q�U��E��H���U��
�E��H���U��J�}� ~�E�P�M��QR�E�P�r�����E��s�}��t!�}��t�M����U���������U���E����E��H�� t9jj j �U�R�o�����E��U�E�#E���u�M��Q�� �E��P���  �e�M����  �U��Bf��+�E�   �M����  f�M�U�R�E�P�M�Q��q�����E�U�;U�t�E��H�� �U��J���  ��E%��  ��]�������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_����������������̋�U��j�hx�h � d�    P���SVW�t�1E�3�P�E�d�    �}�u�����     �x���� 	   ����  �} |�E;��s	�E�   ��E�    �M؉M��}� uhp�j j.h��j証������u̃}� u9�D����     �	���� 	   j j.h��h�hp�����������  �E���M���������D
������؉E�uhċj j/h��j�"�������u̃}� u9�����     ����� 	   j j/h��h�hċ����������   �UR��������E�    �E���M���������D
��t�MQ�n   ���E��4����� 	   �E�����3�uh0�j j9h��j�k�������u��E������   ��MQ�k�����ËE�M�d�    Y_^[��]��̋�U��QV�EP����������t]�}u������   ��u�}u(����HD��tj��������j������;�t�UR�y�����P�!��t	�E�    �	�D �E��EP�`������M���U���������D �}� t�M�Q�C���������3�^��]����̋�U��} uh��j j.hX�j�@�������u̋M�Q��   tK�E�H��t@j�U�BP��C�����M�Q�������E�P�M�    �U�B    �E�@    ]��%� �����̍M��XT���T$�B�J�3��W"������})��������������̍M��(T���T$�B�J�3��'"������M)��������������̋T$�B�J�3���!������%)�������U����   SVW��@����0   ������j �����_^[���   ;������]���U����   SVW��@����0   �����������h��n'����_^[���   ;��K����]�������̋�U��Q3��E���]��U����   SVW��@����0   �����������_^[���   ;�������]�                                                                                                                                                                                                                                                                                                                                    ܥ � � � $� :� N� d� v� �� �� �� �� �� ʦ ަ �� � � .� >� N� \� n� ~� �� �� Ƨ ާ �� � (� 6� D� ^� n� �� �� �� ƨ �  � � 2� >� J� V� h� x� �� �� �� © ̩ ة � �� � � (� >� N� d� t� �� �� �� �� ʪ ت �         � p        �= � p� �� P�        @Z@
��                Data explorer plugin. See the output window ize Cybernetic Genetics data explorer   cg.tiff     c:\program files\maxon\cinema 4d r13\plugins\dataexplorer\cgmenu.cpp    (��   p$ @$ 0# p$ p# �# �# �  �" p$ @$ 0# p$ p# �# �# %s                    �?~   %   res �� (     c:\program files\maxon\cinema 4d r13\resource\_api\c4d_pmain.cpp    ��2     f:\dd\vctools\crt_bld\self_x86\crt\src\dllcrt0.c    @7       �?      �?3      3            �      0C       �       ��              fmod         �; �� /� �� �� �� /� �� -� -� W� -� �� �� /� �� f:\dd\vctools\crt_bld\self_x86\crt\src\onexit.c Unknown Runtime Check Error
   Stack memory around _alloca was corrupted
 A local variable was used before it was initialized
   Stack memory was corrupted
        A cast to a smaller data type has caused a loss of data.  If this was intentional, you should mask the source of the cast with the appropriate bitmask.  For example:  
	char c = (i & 0xFF);
Changing the code in this way will not affect the quality of the resulting optimized code.
    The value of ESP was not properly saved across a function call.  This is usually a result of calling a function declared with one calling convention with a function pointer declared with a different calling convention.
    �%�$t$<$$�#                   Stack around the variable ' ' was corrupted.    The variable '  ' is being used without being initialized.  Run-Time Check Failure #%d - %s Unknown Module Name Unknown Filename        R u n - T i m e   C h e c k   F a i l u r e   # % d   -   % s   R u n t i m e   C h e c k   E r r o r . 
    U n a b l e   t o   d i s p l a y   R T C   M e s s a g e .   Stack corrupted near unknown variable   
   %.2X    Stack around _alloca corrupted  Local variable used before initialization   Stack memory corruption Cast to smaller type causing loss of data   Stack pointer corruption    �(�(�(�(`(        f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ e h \ t y p n a m e . c p p     p N o d e - > _ N e x t   ! =   N U L L     f:\dd\vctools\crt_bld\self_x86\crt\src\tidtable.c   FlsFree FlsSetValue FlsGetValue FlsAlloc    K E R N E L 3 2 . D L L     Client  Ignore  CRT Normal  Free    d*\*X*P*H*Error: memory allocation: bad memory block type.
   Invalid allocation size: %Iu bytes.
    Client hook allocation failure.
    Client hook allocation failure at file %hs line %d.
    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g h e a p . c     _ C r t C h e c k M e m o r y ( )   _ p F i r s t B l o c k   = =   p O l d B l o c k   _ p L a s t B l o c k   = =   p O l d B l o c k     f R e a l l o c   | |   ( ! f R e a l l o c   & &   p N e w B l o c k   = =   p O l d B l o c k )   Error: possible heap corruption at or near 0x%p     p O l d B l o c k - > n L i n e   = =   I G N O R E _ L I N E   & &   p O l d B l o c k - > l R e q u e s t   = =   I G N O R E _ R E Q         _ C r t I s V a l i d H e a p P o i n t e r ( p U s e r D a t a )       The Block at 0x%p was allocated by aligned routines, use _aligned_realloc()     Error: memory allocation: bad memory block type.

Memory allocated at %hs(%d).
 Invalid allocation size: %Iu bytes.

Memory allocated at %hs(%d).
  Client hook re-allocation failure.
 Client hook re-allocation failure at file %hs line %d.
 p U s e r D a t a   ! =   N U L L   _ p F i r s t B l o c k   = =   p H e a d   _ p L a s t B l o c k   = =   p H e a d     p H e a d - > n B l o c k U s e   = =   n B l o c k U s e   p H e a d - > n L i n e   = =   I G N O R E _ L I N E   & &   p H e a d - > l R e q u e s t   = =   I G N O R E _ R E Q         HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.
   HEAP CORRUPTION DETECTED: after %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory after end of heap buffer.

Memory allocated at %hs(%d).
     HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.
       HEAP CORRUPTION DETECTED: before %hs block (#%d) at 0x%p.
CRT detected that the application wrote to memory before start of heap buffer.

Memory allocated at %hs(%d).
 _ B L O C K _ T Y P E _ I S _ V A L I D ( p H e a d - > n B l o c k U s e )     Client hook free failure.
      The Block at 0x%p was allocated by aligned routines, use _aligned_free()    _ m s i z e _ d b g     %hs located at 0x%p is %Iu bytes long.
     %hs located at 0x%p is %Iu bytes long.

Memory allocated at %hs(%d).
   HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.
       HEAP CORRUPTION DETECTED: on top of Free block at 0x%p.
CRT detected that the application wrote to a heap buffer that was freed.

Memory allocated at %hs(%d).
 DAMAGED _heapchk fails with unknown return value!
  _heapchk fails with _HEAPBADPTR.
   _heapchk fails with _HEAPBADEND.
   _heapchk fails with _HEAPBADNODE.
  _heapchk fails with _HEAPBADBEGIN.
 _ C r t S e t D b g F l a g         ( f N e w B i t s = = _ C R T D B G _ R E P O R T _ F L A G )   | |   ( ( f N e w B i t s   &   0 x 0 f f f f   &   ~ ( _ C R T D B G _ A L L O C _ M E M _ D F   |   _ C R T D B G _ D E L A Y _ F R E E _ M E M _ D F   |   _ C R T D B G _ C H E C K _ A L W A Y S _ D F   |   _ C R T D B G _ C H E C K _ C R T _ D F   |   _ C R T D B G _ L E A K _ C H E C K _ D F )   )   = =   0 )     Bad memory block found at 0x%p.
    Bad memory block found at 0x%p.

Memory allocated at %hs(%d).
  _ C r t M e m C h e c k p o i n t   s t a t e   ! =   N U L L   Object dump complete.
  crt block at 0x%p, subtype %x, %Iu bytes long.
 normal block at 0x%p, %Iu bytes long.
  client block at 0x%p, subtype %x, %Iu bytes long.
  {%ld}   %hs(%d) :   #File Error#(%d) :  Dumping objects ->
  Data: <%s> %s
 ( * _ e r r n o ( ) )   _ p r i n t M e m B l o c k D a t a     Detected memory leaks!
 CorExitProcess  m s c o r e e . d l l   f:\dd\vctools\crt_bld\self_x86\crt\src\ioinit.c s t r c p y _ s ( * e n v ,   c c h a r s ,   p )   _ s e t e n v p         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ s t d e n v p . c     f:\dd\vctools\crt_bld\self_x86\crt\src\stdenvp.c    f:\dd\vctools\crt_bld\self_x86\crt\src\stdargv.c    f:\dd\vctools\crt_bld\self_x86\crt\src\a_env.c        �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �      _ c o n t r o l f p _ s ( ( ( v o i d   * ) 0 ) ,   0 x 0 0 0 1 0 0 0 0 ,   0 x 0 0 0 3 0 0 0 0 )   _ s e t d e f a u l t p r e c i s i o n     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i n t e l \ f p 8 . c     s i z e I n B y t e s   >   0   _ c f t o e _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c v t . c     b u f   ! =   N U L L   e+000   s t r c p y _ s ( p ,   ( s i z e I n B y t e s   = =   ( s i z e _ t ) - 1   ?   s i z e I n B y t e s   :   s i z e I n B y t e s   -   ( p   -   b u f ) ) ,   " e + 0 0 0 " )       s i z e I n B y t e s   >   ( s i z e _ t ) ( 3   +   ( n d e c   >   0   ?   n d e c   :   0 )   +   5   +   1 )   _ c f t o e 2 _ l   s i z e I n B y t e s   >   ( s i z e _ t ) ( 1   +   4   +   n d e c   +   6 )     _ c f t o a _ l     _ c f t o f _ l     _ c f t o f 2 _ l   _ c f t o g _ l     ��(�    ( c o u n t   = =   0 )   | |   ( s t r i n g   ! =   N U L L )         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s p r i n t f . c   ( f o r m a t   ! =   N U L L )           �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    pow exp log10   log _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh            �������             ��      �@      �               ���5�h!����?      �?  r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
         R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            �I   hI	   I
   �H   pH   H   �G   pG    G   �F   @F   �E   �E   @E   xD    D!    Bx   �Ay   �Az   �A�   �A�   �AM i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y         w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   e r r o r _ t e x t )     
 
     w c s c a t _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " \ n \ n " )   . . .   w c s n c p y _ s ( p c h ,   p r o g n a m e _ s i z e   -   ( p c h   -   p r o g n a m e ) ,   L " . . . " ,   3 )   < p r o g r a m   n a m e   u n k n o w n >     w c s c p y _ s ( p r o g n a m e ,   p r o g n a m e _ s i z e ,   L " < p r o g r a m   n a m e   u n k n o w n > " )     R u n t i m e   E r r o r ! 
 
 P r o g r a m :     w c s c p y _ s ( o u t m s g ,   ( s i z e o f ( o u t m s g )   /   s i z e o f ( o u t m s g [ 0 ] ) ) ,   L " R u n t i m e   E r r o r ! \ n \ n P r o g r a m :   " )     _ N M S G _ W R I T E   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c r t 0 m s g . c     M S P D B 1 0 0 . D L L     r   PDBOpenValidate5    E n v i r o n m e n t D i r e c t o r y         S O F T W A R E \ M i c r o s o f t \ V i s u a l S t u d i o \ 1 0 . 0 \ S e t u p \ V S   RegCloseKey RegQueryValueExW    RegOpenKeyExW   A D V A P I 3 2 . D L L     ... Assertion Failed    Error   Warning �O�O�O    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t . c   Microsoft Visual C++ Debug Library  _CrtDbgReport: String too long or IO Error  s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )     Debug %s!

Program: %s%s%s%s%s%s%s%s%s%s%s%s

(Press Retry to debug the application)    
Module:    
File:  
Line:  

  Expression:     

For information on how your program can cause an assertion
failure, see the Visual C++ documentation on asserts.      m e m c p y _ s ( s z S h o r t P r o g N a m e ,   s i z e o f ( T C H A R )   *   ( 2 6 0   -   ( s z S h o r t P r o g N a m e   -   s z E x e N a m e ) ) ,   d o t d o t d o t ,   s i z e o f ( T C H A R )   *   3 )     <program name unknown>  s t r c p y _ s ( s z E x e N a m e ,   2 6 0 ,   " < p r o g r a m   n a m e   u n k n o w n > " )     _ _ c r t M e s s a g e W i n d o w A   A s s e r t i o n   F a i l e d     E r r o r   W a r n i n g    T�S�S    M i c r o s o f t   V i s u a l   C + +   D e b u g   L i b r a r y     _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r     w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )   D e b u g   % s ! 
 
 P r o g r a m :   % s % s % s % s % s % s % s % s % s % s % s % s 
 
 ( P r e s s   R e t r y   t o   d e b u g   t h e   a p p l i c a t i o n )     
 M o d u l e :     
 F i l e :     
 L i n e :     E x p r e s s i o n :           
 
 F o r   i n f o r m a t i o n   o n   h o w   y o u r   p r o g r a m   c a n   c a u s e   a n   a s s e r t i o n 
 f a i l u r e ,   s e e   t h e   V i s u a l   C + +   d o c u m e n t a t i o n   o n   a s s e r t s .     w c s c p y _ s ( s z E x e N a m e ,   2 6 0 ,   L " < p r o g r a m   n a m e   u n k n o w n > " )   _ _ c r t M e s s a g e W i n d o w W   f:\dd\vctools\crt_bld\self_x86\crt\src\mlock.c  ( L " B u f f e r   i s   t o o   s m a l l "   & &   0 )   B u f f e r   i s   t o o   s m a l l   ( ( ( _ S r c ) ) )   ! =   N U L L     s t r c p y _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c p y _ s . i n l   ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n B y t e s ) )   >   0      Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(    �^�^�^�^�^�^�^�^�^�^�^ )x^p^l^h^d^`^\^X^T^H^D^@^<^8^4^0^,^(^$^�" ^^^^^^�"^^ ^�]�]�]�]�]�]�]�]�]�]�]�]�]�]�]�]�]p]P]0]]�\�\�\�\l\L\$\\�[�[�[�[�[�[�[�[x[X[0[[�Z�Z�ZtZPZ$Z�Y�Y )�Y�Y�YxY\Y    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l o c a l r e f . c       ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   ! =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   ! =   N U L L ) )   | |   ( ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w l o c a l e   = =   N U L L )   & &   ( p t l o c i - > l c _ c a t e g o r y [ c a t e g o r y ] . w r e f c o u n t   = =   N U L L ) )     H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun f:\dd\vctools\crt_bld\self_x86\crt\src\mbctype.c    _ e x p a n d _ b a s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e x p a n d . c   p B l o c k   ! =   N U L L     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s c t y p e . c     ( u n s i g n e d ) ( c   +   1 )   < =   2 5 6     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w i n s i g . c   ( " I n v a l i d   s i g n a l   o r   e r r o r " ,   0 )     r a i s e   _ c o n t r o l f p _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ t r a n \ c o n t r l f p . c   ( " I n v a l i d   i n p u t   v a l u e " ,   0 )     p f l t   ! =   N U L L         s i z e I n B y t e s   >   ( s i z e _ t ) ( ( d i g i t s   >   0   ?   d i g i t s   :   0 )   +   1 )   _ f p t o s t r     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f p t o s t r . c       s t r c p y _ s ( r e s u l t s t r ,   r e s u l t s i z e ,   a u t o f o s . m a n )     _ f l t o u t 2     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ c f o u t . c         ( " i n c o n s i s t e n t   I O B   f i e l d s " ,   s t r e a m - > _ p t r   -   s t r e a m - > _ b a s e   > =   0 )     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f l s b u f . c     s t r   ! =   N U L L   ( n u l l )     (null)             EEE50 P    ( 8PX 700WP        `h````  xpxxxx          f:\dd\vctools\crt_bld\self_x86\crt\src\output.c     ( " ' n '   f o r m a t   s p e c i f i e r   d i s a b l e d " ,   0 )     ( c h   ! =   _ T ( ' \ 0 ' ) )     (   ( _ S t r e a m - > _ f l a g   &   _ I O S T R G )   | |   (   f n   =   _ f i l e n o ( _ S t r e a m ) ,   (   ( _ t e x t m o d e _ s a f e ( f n )   = =   _ _ I O I N F O _ T M _ A N S I )   & &   ! _ t m _ u n i c o d e _ s a f e ( f n ) ) ) )   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o u t p u t . c   ( s t r e a m   ! =   N U L L )     _ s e t _ e r r o r _ m o d e       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ e r r m o d e . c     ( " I n v a l i d   e r r o r _ m o d e " ,   0 )   GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L         ( L " S t r i n g   i s   n o t   n u l l   t e r m i n a t e d "   & &   0 )   S t r i n g   i s   n o t   n u l l   t e r m i n a t e d   w c s c a t _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s c a t _ s . i n l   ( ( _ D s t ) )   ! =   N U L L   & &   ( ( _ S i z e I n W o r d s ) )   >   0     w c s n c p y _ s   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ t c s n c p y _ s . i n l     w c s c p y _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m a l l o c . h   ( " C o r r u p t e d   p o i n t e r   p a s s e d   t o   _ f r e e a " ,   0 )       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ d b g r p t t . c         _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g     w c s c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )         e   =   m b s t o w c s _ s ( & r e t ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )       s t r c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )   %s(%d) : %s     s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ n " )          s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   " \ r " )   s t r c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )         s t r c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   " A s s e r t i o n   f a i l e d :   "   :   " A s s e r t i o n   f a i l e d ! " )     Assertion failed!   Assertion failed:       s t r c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )   , Line  <file unknown>  Second Chance Assertion Failed: File    _ i t o a _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )   _ V C r t D b g R e p o r t A   w c s t o m b s _ s ( & r e t ,   s z a O u t M e s s a g e ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )   _CrtDbgReport: String too long or Invalid characters in String      s t r c p y _ s ( s z O u t M e s s a g e 2 ,   4 0 9 6 ,   " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I n v a l i d   c h a r a c t e r s   i n   S t r i n g " )   w c s t o m b s _ s ( ( ( v o i d   * ) 0 ) ,   s z O u t M e s s a g e 2 ,   4 0 9 6 ,   s z O u t M e s s a g e ,   ( ( s i z e _ t ) - 1 ) )         w c s c p y _ s ( s z O u t M e s s a g e ,   4 0 9 6 ,   s z L i n e M e s s a g e )   % s ( % d )   :   % s   w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ n " )        w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   L " \ r " )         w c s c a t _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z U s e r M e s s a g e )         w c s c p y _ s ( s z L i n e M e s s a g e ,   4 0 9 6 ,   s z F o r m a t   ?   L " A s s e r t i o n   f a i l e d :   "   :   L " A s s e r t i o n   f a i l e d ! " )     A s s e r t i o n   f a i l e d !   A s s e r t i o n   f a i l e d :           w c s c p y _ s ( s z U s e r M e s s a g e ,   4 0 9 6 ,   L " _ C r t D b g R e p o r t :   S t r i n g   t o o   l o n g   o r   I O   E r r o r " )     
   ,   L i n e     < f i l e   u n k n o w n >     S e c o n d   C h a n c e   A s s e r t i o n   F a i l e d :   F i l e         _ i t o w _ s ( n L i n e ,   s z L i n e M e s s a g e ,   4 0 9 6 ,   1 0 )   _ V C r t D b g R e p o r t W   GetUserObjectInformationA   MessageBoxA s i z e I n B y t e s   > =   c o u n t     s r c   ! =   N U L L   m e m c p y _ s     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m e m c p y _ s . c   d s t   ! =   N U L L                                                                                                                                                                                                                                                                                         ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������_ v s n p r i n t f _ h e l p e r   ( " B u f f e r   t o o   s m a l l " ,   0 )       s t r i n g   ! =   N U L L   & &   s i z e I n B y t e s   >   0   _ v s p r i n t f _ s _ l   f o r m a t   ! =   N U L L     _ v s n p r i n t f _ s _ l     	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~  _ _ s t r g t o l d 1 2 _ l         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ i n c l u d e \ s t r g t o l d 1 2 . i n l     _ L o c a l e   ! =   N U L L   1#QNAN  s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # Q N A N " )     1#INF   s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N F " )   1#IND       s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # I N D " )   1#SNAN      s t r c p y _ s ( f o s - > m a n ,   2 1 + 1 ,   " 1 # S N A N " )     $ I 1 0 _ O U T P U T   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ p r e b u i l d \ c o n v \ x 1 0 f o u t . c     ( " I n v a l i d   f i l e   d e s c r i p t o r .   F i l e   p o s s i b l y   c l o s e d   b y   a   d i f f e r e n t   t h r e a d " , 0 )   ( _ o s f i l e ( f h )   &   F O P E N )   _ l s e e k i 6 4       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ l s e e k i 6 4 . c       ( f h   > =   0   & &   ( u n s i g n e d ) f h   <   ( u n s i g n e d ) _ n h a n d l e )     _ w r i t e     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w r i t e . c     i s l e a d b y t e ( _ d b c s B u f f e r ( f h ) )   ( ( c n t   &   1 )   = =   0 )     _ w r i t e _ n o l o c k   ( b u f   ! =   N U L L )   f:\dd\vctools\crt_bld\self_x86\crt\src\_getbuf.c    f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ g e t b u f . c     _ i s a t t y       f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ i s a t t y . c   f:\dd\vctools\crt_bld\self_x86\crt\src\_file.c  _ f i l e n o   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f i l e n o . c   _ w c t o m b _ s _ l   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c t o m b . c   s i z e I n B y t e s   < =   I N T _ M A X     _ m b s t o w c s _ l _ h e l p e r     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b s t o w c s . c   s   ! =   N U L L   r e t s i z e   < =   s i z e I n W o r d s     b u f f e r S i z e   < =   I N T _ M A X   _ m b s t o w c s _ s _ l   ( p w c s   = =   N U L L   & &   s i z e I n W o r d s   = =   0 )   | |   ( p w c s   ! =   N U L L   & &   s i z e I n W o r d s   >   0 )   s t r c a t _ s     l e n g t h   <   s i z e I n T C h a r s   2   < =   r a d i x   & &   r a d i x   < =   3 6       s i z e I n T C h a r s   >   ( s i z e _ t ) ( i s _ n e g   ?   2   :   1 )   s i z e I n T C h a r s   >   0     x t o a _ s         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ x t o a . c   _ w c s t o m b s _ l _ h e l p e r         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ w c s t o m b s . c   p w c s   ! =   N U L L     s i z e I n B y t e s   >   r e t s i z e   _ w c s t o m b s _ s _ l   ( d s t   ! =   N U L L   & &   s i z e I n B y t e s   >   0 )   | |   ( d s t   = =   N U L L   & &   s i z e I n B y t e s   = =   0 )   _ v s w p r i n t f _ h e l p e r   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ v s w p r i n t . c       s t r i n g   ! =   N U L L   & &   s i z e I n W o r d s   >   0   _ v s n w p r i n t f _ s _ l   x t o w _ s     ��bad exception   T���0	    ( ( s t a t e   = =   S T _ N O R M A L )   | |   ( s t a t e   = =   S T _ T Y P E ) )         ( " I n c o r r e c t   f o r m a t   s p e c i f i e r " ,   0 )       ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp       _ o u t p u t _ s _ l   _ g e t _ o s f h a n d l e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ o s f i n f o . c         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ m b t o w c . c   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   1   | |   _ l o c _ u p d a t e . G e t L o c a l e T ( ) - > l o c i n f o - > m b _ c u r _ m a x   = =   2     _ w o u t p u t _ s _ l     ( s t r   ! =   N U L L )   csm�               �        ԝ0	Unknown exception   C O N O U T $   f c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ f c l o s e . c   _ f c l o s e _ n o l o c k     ( _ o s f i l e ( f i l e d e s )   &   F O P E N )     _ c o m m i t   f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c o m m i t . c   ( f i l e d e s   > =   0   & &   ( u n s i g n e d ) f i l e d e s   <   ( u n s i g n e d ) _ n h a n d l e )     _ c l o s e         f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ c l o s e . c     f : \ d d \ v c t o o l s \ c r t _ b l d \ s e l f _ x 8 6 \ c r t \ s r c \ _ f r e e b u f . c   s t r e a m   ! =   N U L L         H                                                           t��               �<�           L�\�x���    �       ����    @   <��       ����    @   ��           ��x���    8�        ����    @   ̜           ܜ��                ���            8�̜            T� �           0�8�    T�        ����    @    �            ؿh�           x�����    ؿ       ����    @   h���        ����    @   ��           ̝��                ����         �  ��  �? �@  C h � �     P2         �2     ����    ����    ����    g4     ����    ����    �����6  7     ����    ����    ����    K<     ����    ����    ����$A *A     ����    ����    �����A �A     ����    ����    ����    +D     ����    ����    ����    �H ����    �H ����    ����    ����    hK ����    �K ����    ����    ����    <Q     ����    ����    ����    �R     ����    ����    ����    AY     ����    ����    ����    `     ����    ����    ����    �d     ����    ����    ����    �e     ����    ����    ����    {h     ����    ����    ����    �l     ����    ����    ����    �s     ����    ����    ������ '�     ����    ����    ����    �     ����    ����    ����    ��     ����    ����    ����    ��     ����    ����    ����    n� ����`"�   ��                       ����    ����    ������ ��     ����    ����    ������ ��     ����    ����    ����=� C�     ����    ����    ����    �����"�   ��                       ����    ����    ����    �/        u.����    |��    ����    9        �6����    ����    ����    �Z    ����    ����    ����    $�    ����    ����    ����    ?�    ��    ��   ����    ؿ    ����       ��    ��    ����       �����    ����    ����    ��    ��������    ����    ����    ��    ��������    ����    ����F�L�    ����    ����    ����U�[�    ����    ����    ������@           ������    ����                  t�"�   ��   ��                   ����    ����    ����    ��    ����    ����    ����    �    ����    ����    ����    ��        ������    ����    ����    Q    ����    ����    ����    u    ����    ����    ����    ���         ��                        ܥ � � � $� :� N� d� v� �� �� �� �� �� ʦ ަ �� � � .� >� N� \� n� ~� �� �� Ƨ ާ �� � (� 6� D� ^� n� �� �� �� ƨ �  � � 2� >� J� V� h� x� �� �� �� © ̩ ة � �� � � (� >� N� d� t� �� �� �� �� ʪ ت �     �GetCurrentThreadId  � DecodePointer �GetCommandLineA � EncodePointer WideCharToMultiByte  IsDebuggerPresent gMultiByteToWideChar �RaiseException  EGetProcAddress  ?LoadLibraryW  �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree GetModuleHandleW  �InterlockedIncrement  sSetLastError  GetLastError  �InterlockedDecrement  �HeapValidate  �IsBadReadPtr  ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter IsProcessorFeaturePresent GetModuleFileNameW  %WriteFile �HeapFree  �HeapAlloc JGetProcessHeap  �VirtualQuery  bFreeLibrary � EnterCriticalSection  9LeaveCriticalSection  RtlUnwind hGetACP  7GetOEMCP  rGetCPInfo 
IsValidCodePage �HeapReAlloc �HeapSize  �HeapQueryInformation  �OutputDebugStringA  $WriteConsoleW �OutputDebugStringW  -LCMapStringW  iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll              нQ    B�          8� <� @� �)  S�   dataexplorer.dll c4d_main                                                                                                                                                                        �"    .?AVCGMenu@@    �"    .?AVCommandData@@   �"    .?AVBaseData@@  Q   �"    .?AVtype_info@@ u�  s�  N�@���D                               ��������   ����   ��������    �����
                                                          0000000000?         �@   �@   �@   �@   0A   (A!    A   �@   �@   �@   A   A   p@   l@    h@   �@   |@   A   t@    A   �@   �@   �@   �@"   �@#   �@$   �@%   �@&   �@      �      ���������              �       �D        � 0            �O0L                                                                                                                                                                                                                                                                                     C       �e�e�e�e�e�e�e�e�e�e�e�e�e|exetepelehede`e\eXeTePeLeDe8e0e(ehe eeee�d�d�d�d�d�d�d�d	         �d�d�d�d�d�dxdhdXdHd4d dd�c�c�c�c�c�c�c�c�c�c�c�c�c�cxclc`c�cTcHc8c$cc c�b�b�b�b�b�b                                                                                           ��            ��            ��            ��            ��                              ȼ        ������ �                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��                                     	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 `� ����        �k�k�&  ����         ������������         �            .   .   ��H�H�H�H�H�H�H�H�H�ļL�L�L�L�L�L�L�ȼ���   ���5      @   �  �   ����             ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �"    .?AVbad_exception@std@@ �"    .?AVexception@std@@                .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
    ����                                                                                                                                                                                                                                                                                               �                 0  �              	  H   X� Z  �      <assembly xmlns="urn:schemas-microsoft-com:asm.v1" manifestVersion="1.0">
  <trustInfo xmlns="urn:schemas-microsoft-com:asm.v3">
    <security>
      <requestedPrivileges>
        <requestedExecutionLevel level="asInvoker" uiAccess="false"></requestedExecutionLevel>
      </requestedPrivileges>
    </security>
  </trustInfo>
</assembly>PAPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPADDINGPADDINGXXPAD   h   &0�0�0�01B1�12_2d2m2�2�2�2�3�4c6�6#7E7�7�7;8�89=9�9:�:�:�:�:;*;�;k<�<=�=�=�=�=�=�=;>�?�?�?    l   0�0�0�15555$5+52595@5h5�5�5�6�67`7�78�8�9�9�9:::R:W:`:�:�:�:�:�:;;U;|;�;�;�;�;�;<�=?�? 0  �   0h0�0R2e2�283=3O3�3�3�3444(414>4o4�4�4�4�4�4�5�5�5�5�5�5y6�6�6�6g7k7q7u7{77�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7*8C8�8�8�8�89.9�9M:�;�;�;�;<y<�<�<�<=9=z==�=�=�=�=>>>>P>W>r>�>�>B?f?�?�? @  T  000a0�0�0�0�01X1]1o1�1�12R2�2�2�2�2�233!363H3M3_3�3�3�3�35'575>5M5T5`5g5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�56666"6(6.646:6?6D6J6O6U6^6e6l6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67/767=7`7�7�7�7�7�7�7�7�7�7�7�7�788&8b8�8�89"9?9c9i9p9�9�9:::�:;;F;�;�;<%<,<6<=<D<P<W<^<o<y<�<�<�=�=�=�=�=>> >6>B>K>P>Y>e>n>�>�>�>�>�>?k?p?�?�?   P  @  0*030;0D0L0R0X0`0f0l0t0�0�0�0�0�01�1H2M2_2?3H3Q3a3m3�3�3�3�3�3�3�3�3�344U4v4�4�4�4555r5~5�5�56!6�6�6�6�6�6�6�6�6�6�67
7777&7,7Q7m7�7�788&8B8`8j8v8�8�8�8�8�8�8�8�8�8h9p9y9�9�9�9�9�9�9�9&:A:M:R:�:�:�:�:;;d;j;�;�;�;<$<\<b<�<�<�<==1=:=?=e=o={=�=�=�=�=�=�='>H>M>_>�>�>�>�>�>�>�>�> ??"?.?7?]?i?�?�?   `  �   x0}0�0�0111,111N1S1p1u1�1�1�1*262?2�2�2�23N3�3�3�324a4�4�4�4�4�4�4�45;5G5t5y5~5�5�5�5�5�5�5e6l6�6�6�6�6�6�677.7k7878[8f8)9:9R9c9:::K:P:y:�:
;;E;g;�;�;�;�;1<�<�<�<=><>A>F>~>�>?,?1?w?�?�?�?�?�?�?�?   p  �    000030�0�0�01;1J1U1f1w1~1�1�1�1�1�1�1�1�1�1�1�1�1222@2M2Y2i2p2�2�2�23333Q3V3c3h3v3�3�3�3�344G4n5x5�5�5�5�6�6�6�6�6�6�6�7�7�7C8�8�89^9e9�9�9�9�9�9�9:.:|:�:�:�:�:;);>;C;H;|;�;�;�;�;�;�;�;�;�;
<<e<�<�<�<   �  �   Q0�0�0�0
1-1D1K1^1t1{1�1�1�1�1�1�1�1-2�2�23/3}384C4P4X4g4|4�4�4�4�4�4�5�5�5Q7d7�7�7�7�:�:�:;";';L;X;�;�;�;~<�<�<�<�<�<�<,=1=6=x=�=�=�=�=�>�>�>�>�? �  x   �0�0�0�0�01#1P1U1Z1�1�1�1�1�18d8p8�8�8�8�8�89
99�9�9,:1:6:h:t:�:�:�:)<x<�<�<�<�<�<�<==#=�?�?�?�?�?�?�?�?�? �  �   00000$0+030;0C0O0X0]0c0m0w0�0�0�0�0�0�0�0�0�0�0�1�1�1�12272E2�2�2)3u3�3�34d4�4�495T5�5�5=6�6�6�6�6A7L7�7�7�78U8`8�8�89Y9�9�9J:�:�:�: ;;;;;;;; ;$;(;,;0;4;�;�;�;�;�;�;�;�; <<<<<<><�<y=~=W>�>-? �  P   S3�3�4�4�4�4�5�56"6E6P6s6~67$9392<G<\<�<�<�<�<�<,=�=�=5>�>�>�>�>??   �  �   0�0(1�1�1�1D2�2�2�2y3�344)4P4U4Z4_4i4�4�4�4�4�45"5'5.5i5n5s5x5�5�5�5�5�5�5�5	676T6�6�6�6�6�6�6�6578
8�8�8�8�89999:9?9b9p9�9�9�9�9X:^:m:v::�:�:�:@;~;�;�;�;�;�;�; <<�<�<�<�<�<�<�<="=.=I=Y=e=�=�=�=�=�=0>6>d>i>n>�>�>�>�>�>�?�?   �  �    00
00h0m0r0y0�01&1@1L1`1l1�1�1�1�1�1�12"2.2>2J2�2�2�2�2�233 3%3L3�3�3�3�344V4c4p4}4�4�4�4�4�4�4�45+5T5k5�5�5�5K6r6y6�6�6�6�67	77Q7Y7�7�7�7�7�7U8]8�8�8�8�8�8�8.959<:�:�:�:;%;4;Y;g;t;�;�;�;�<�<=U=a=l>�>�>�> ??E?k?�?�?�?�?   �  �   0*0F0o0�0�0�01g2�2O3[3-4X4]4o4�4�4(5-5?5b5�5�5�5�5�5�586=6O6�67797N7t77�7�7�78"8)83878@8R8\8�8�8�89#9-9R9\9�9�9?:�:�:Y;�;�;�<T=[=�=�=�=�=�=H>w>�>�>   �  �   �1�1W2c2�2�23'3.3w3�3�3�3�3�3%4,4>4E4v4�4�4U5\5�5�5�56	6�6�6�6�6�8�899#9(9,909Y99�9�9�9�9�9�9�9�9�9
:::::�:�:�:�:�:�:�:�:;9;@;D;H;L;P;T;X;\;�;�;�;�;�;�<�<=(=>>!>8>=>O>�>�>�>??y?�?�?�?�?�?�?   �   000:0W0t0�0�0&1+101J1�1�1�1�2�2�2�2�2�2�2�2&3-3I3x3�3�4�4�4�4�4�5�7	89J:S:}:�:�:�:�:�:�:�:$;-;W;\;a;�;�;�;�;�;�<8===B=
?<?T?[?c?h?l?p?�?�?�?�?�?�?�?�?�?�?        0J0P0T0X0\0�0�0�0�0�0�0�01G1y1�1�1�1�1�1�1�1�1�1�1�1�1�1_4h4�5�5f6r6�7�7�8094989<9@9D9H9L9{9�9�9�9�9�9�9�9:H:T:Z:o:y:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;;;;$;.;5;>;E;�;�;�;�;�;�;�;�;a<j<�<�<�<�<�<*=3=]=b=g=�=�=>:>C>m>r>w>�>�>%?N?W?�?�?�?�?�?       j0s0�0�0�0�0�0R1Y1�1�1�1�1�1F2O2�2323[3d3�3�3�3�3�3�4�4�4�4�455Z5c5�5�5�56$6Q6z6�6�6�6�6�6�6�7�7�7�78�8�8�8�89+919L9Y9^9d9q9v9|9�9�9:8:=:B:G:z:�:�:�:�:�:�:�:
;; ;%;*;S;X;];b;�;�;�;�;3<8<=<B<m<r<w<�<�<�<==!=&=I=R=�=�=�>�>�>�>$?+?5?G?Q?o?t?y?�?�?   0 (  (0-0F011-12171_1e1�1�1�1�1�1�1�1"2'2,2b2g2l2q2�2�2�2�2�2�2�2 343E3J3O3T3}3�3�3�3�34"4'4]4b4g4l4�4�4�4�4�4�4,51565;5^5g5�56�6�6�67!7(7c7j7y7�7�7�788Z8a8k8}8�8�8�8�89$9Y9�9�9�9�9�9�9�9�9�9�9�9�9:	::::*:/:5:=:G:N:S:Y:d:n:u:~:�:�:�:�:;;;5;<;�;�;�;�;�;"<+<U<Z<_<�<�<�<�<�<�>R?W? @ L   00050�2Q3]3�3�3�3�:�:�:;";X;w;�;�;�;�;<1<P<o<�<�<�<�=U>}>�>[?�?�? P �   �0`11�1�1222Y2b2�2�2�2�3�3�3�3�324>4k4p4u4�4�4�4/5;5h5m5r5�5�5)656b6g6l6�6�6�6 77G7�7�7�7i8q8�8�8�8 99B9J9H:M:_:t:x:�:�:�:P<o<x<   ` (   v2�29<9�9�9�9�9�9�:�;�;==>> p `   �2�2�2�2�2�2�2�2�2�2�2 33333P3T3X3�3�3�3�3�34�4�9�:�:�:�:@;E;J;O;�;�;�;�;�;�;�;�;   � �   000r0�0�0�0�0�011'1\1a1f1�1�12�2�2�2�23&3H3M3_3�3�3�344424J4S4�4�4�4�455�5�5�566626f6o6�6�6�6�67W7a7�7�7 88#8I8n8�89�9�9�9:U:_:�:�:;D;d<n<�<�=�=�=??e?o?�?�?�? � �   0`0�0�0�0�0�0�1�1�1222-2F2X2a2m2v2�2�2�2�2�2�2�2�2�233B3^3z3�3�3�3�3�3�34g4x4�4�4�45)525\5a5f5�5�5�56/64696�6�6777�7�78858:8?8)929\9a9f9*:R:B;�;t<�<�<�<�<�< =v=�=�=�=�=->4>�>�>??F?K?P? � �   00D0I0N0�0�0�0�0	111�1�1�1�1�1222�2�2�2�2�2"3'3,3l3t3;4D4n4s4x4�4�4�4�4�455^5g5�5�5�5�5�5666�6�677$7�7�7�7	888<9�9�9g:<= =M=R=W=�=�=>>?>D>I>�>�>3?:?t?�?�?�?�?   � �   o0{0�0�0�0�0�0(1-121�2�2�2�2�2R3^3�3�3�3�344�455^5j5�5�5�5�5�5�6�67#7(7M7V7�7�7�7�7�788E8J8O8�8�8�8�8�8�9�9�9�9�9P=]= � <   j0�0�0�3�3�3666999x;};�;�<�<�<H>X>�>�>|?�?�?   � p   !0&0+0�0�011Z1f1�1�1�1�1�12#2(2�23N3Z3�3�3�3�3P4\4�4�4�4@5G5U6\6�7�7n899�9F:R:�:�:�:g;�;�;< <O<V<   � �   �1�1!2&2+2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�233333 3$3(3,3034383<3@3D3�57!7E7Q7x7�7�7�78:8F8~8�8�8�8�8�8
99979X9]9o9�9�9":-:g:r:�:�:�:�:=;F;<�<==/=q==�=�=�=�=�=�=�?�?�?�?�? � h   	0#0C0_0�0�0�0<1�1�1�1�1�1-292i2n2s23Q3�3�3�3�3�3,4�4�4�5�5	77�7�899�9�9%:*:/:;�;�;�;�;�;�;     �   �1�1�1�1�12 2$2(2,2024282<2@2D2H2L2P2h2l2p2t2x2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2Y4�4�4$505�56�7�7N8�89R9%:+:0:G:P:X:_:x:}:�:�:�:�:�:�:�;�;�;�;�;�<�<�<�<�<=,=1=6=\=t=}=�=�=�=�=>>J>S>�>�>  T   10=0�0�0�1�12Q2t2}2�2�2�2�2�2383=3B3{3�3�3 474m4�4�4�4�4V5z5�5�56?6I6�6     �   $1(1,181<1@1D1H1T1X1\122 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2�2�2�2�23�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�6�6�6�6�6�699999l:p:t:x:|: 0    $?(? @ <   $:,:4:<:D:L:T:\:d:l:t:|:�:�:�:�:�:�:�:�:�:�:�?�?�?   P �   444�>�> ???????? ?$?(?,?0?4?8?<?@?D?H?L?P?T?X?\?`?d?h?l?p?t?x?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   ` H    00000000 0$0(0,0004080<0@0D0H0L0P0T0X0\0`0d0h0l0p0t0x0   � �   �5�5�5�5999< <4<8<H<L<P<T<\<t<x<�<�<�<�<�<�<�<�<�<�<====,=0=8=P=`=d=t=x=|=�=�=�=�=�=�=�=�=> >@>\>`>�>�>�>�>�>�> ??(?4?P?p?�?�?�?�? � |   000P0l0p0�0�0�0�0�014181T1X1t1x1�1�1�1�1�12202P2p2x2�2�2�2�2�2�2�2�2�2�2333,303L3P3l3p3�3�3�3�3�34(444P4p4�4 � `  0080T0 11111111 1$141<1D1L1T1\1d1l1t1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1222d2h2�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,4044484<4@4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4X5h5x5�5�5�5�5�5�5�5�5:p<�<�<�<�<�<�<�<�<�<�<�<�<�<�< ======== =$=X=`=�?�?                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    